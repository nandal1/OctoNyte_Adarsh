module RegFileMT2R1WVec (
	clock,
	reset,
	io_threadID,
	io_src1,
	io_src2,
	io_dst1,
	io_wen,
	io_dst1data,
	io_src1data,
	io_src2data
);
	input clock;
	input reset;
	input [1:0] io_threadID;
	input [4:0] io_src1;
	input [4:0] io_src2;
	input [4:0] io_dst1;
	input io_wen;
	input [31:0] io_dst1data;
	output wire [31:0] io_src1data;
	output wire [31:0] io_src2data;
	wire [1:0] io_threadID_0 = io_threadID;
	wire [4:0] io_src1_0 = io_src1;
	wire [4:0] io_src2_0 = io_src2;
	wire [4:0] io_dst1_0 = io_dst1;
	wire io_wen_0 = io_wen;
	wire [31:0] io_dst1data_0 = io_dst1data;
	wire [31:0] _regs_WIRE_0 = 32'h00000000;
	wire [31:0] _regs_WIRE_1 = 32'h00000000;
	wire [31:0] _regs_WIRE_2 = 32'h00000000;
	wire [31:0] _regs_WIRE_3 = 32'h00000000;
	wire [31:0] _regs_WIRE_4 = 32'h00000000;
	wire [31:0] _regs_WIRE_5 = 32'h00000000;
	wire [31:0] _regs_WIRE_6 = 32'h00000000;
	wire [31:0] _regs_WIRE_7 = 32'h00000000;
	wire [31:0] _regs_WIRE_8 = 32'h00000000;
	wire [31:0] _regs_WIRE_9 = 32'h00000000;
	wire [31:0] _regs_WIRE_10 = 32'h00000000;
	wire [31:0] _regs_WIRE_11 = 32'h00000000;
	wire [31:0] _regs_WIRE_12 = 32'h00000000;
	wire [31:0] _regs_WIRE_13 = 32'h00000000;
	wire [31:0] _regs_WIRE_14 = 32'h00000000;
	wire [31:0] _regs_WIRE_15 = 32'h00000000;
	wire [31:0] _regs_WIRE_16 = 32'h00000000;
	wire [31:0] _regs_WIRE_17 = 32'h00000000;
	wire [31:0] _regs_WIRE_18 = 32'h00000000;
	wire [31:0] _regs_WIRE_19 = 32'h00000000;
	wire [31:0] _regs_WIRE_20 = 32'h00000000;
	wire [31:0] _regs_WIRE_21 = 32'h00000000;
	wire [31:0] _regs_WIRE_22 = 32'h00000000;
	wire [31:0] _regs_WIRE_23 = 32'h00000000;
	wire [31:0] _regs_WIRE_24 = 32'h00000000;
	wire [31:0] _regs_WIRE_25 = 32'h00000000;
	wire [31:0] _regs_WIRE_26 = 32'h00000000;
	wire [31:0] _regs_WIRE_27 = 32'h00000000;
	wire [31:0] _regs_WIRE_28 = 32'h00000000;
	wire [31:0] _regs_WIRE_29 = 32'h00000000;
	wire [31:0] _regs_WIRE_30 = 32'h00000000;
	wire [31:0] _regs_WIRE_31 = 32'h00000000;
	wire [31:0] _regs_WIRE_32 = 32'h00000000;
	wire [31:0] _regs_WIRE_33 = 32'h00000000;
	wire [31:0] _regs_WIRE_34 = 32'h00000000;
	wire [31:0] _regs_WIRE_35 = 32'h00000000;
	wire [31:0] _regs_WIRE_36 = 32'h00000000;
	wire [31:0] _regs_WIRE_37 = 32'h00000000;
	wire [31:0] _regs_WIRE_38 = 32'h00000000;
	wire [31:0] _regs_WIRE_39 = 32'h00000000;
	wire [31:0] _regs_WIRE_40 = 32'h00000000;
	wire [31:0] _regs_WIRE_41 = 32'h00000000;
	wire [31:0] _regs_WIRE_42 = 32'h00000000;
	wire [31:0] _regs_WIRE_43 = 32'h00000000;
	wire [31:0] _regs_WIRE_44 = 32'h00000000;
	wire [31:0] _regs_WIRE_45 = 32'h00000000;
	wire [31:0] _regs_WIRE_46 = 32'h00000000;
	wire [31:0] _regs_WIRE_47 = 32'h00000000;
	wire [31:0] _regs_WIRE_48 = 32'h00000000;
	wire [31:0] _regs_WIRE_49 = 32'h00000000;
	wire [31:0] _regs_WIRE_50 = 32'h00000000;
	wire [31:0] _regs_WIRE_51 = 32'h00000000;
	wire [31:0] _regs_WIRE_52 = 32'h00000000;
	wire [31:0] _regs_WIRE_53 = 32'h00000000;
	wire [31:0] _regs_WIRE_54 = 32'h00000000;
	wire [31:0] _regs_WIRE_55 = 32'h00000000;
	wire [31:0] _regs_WIRE_56 = 32'h00000000;
	wire [31:0] _regs_WIRE_57 = 32'h00000000;
	wire [31:0] _regs_WIRE_58 = 32'h00000000;
	wire [31:0] _regs_WIRE_59 = 32'h00000000;
	wire [31:0] _regs_WIRE_60 = 32'h00000000;
	wire [31:0] _regs_WIRE_61 = 32'h00000000;
	wire [31:0] _regs_WIRE_62 = 32'h00000000;
	wire [31:0] _regs_WIRE_63 = 32'h00000000;
	wire [31:0] _regs_WIRE_64 = 32'h00000000;
	wire [31:0] _regs_WIRE_65 = 32'h00000000;
	wire [31:0] _regs_WIRE_66 = 32'h00000000;
	wire [31:0] _regs_WIRE_67 = 32'h00000000;
	wire [31:0] _regs_WIRE_68 = 32'h00000000;
	wire [31:0] _regs_WIRE_69 = 32'h00000000;
	wire [31:0] _regs_WIRE_70 = 32'h00000000;
	wire [31:0] _regs_WIRE_71 = 32'h00000000;
	wire [31:0] _regs_WIRE_72 = 32'h00000000;
	wire [31:0] _regs_WIRE_73 = 32'h00000000;
	wire [31:0] _regs_WIRE_74 = 32'h00000000;
	wire [31:0] _regs_WIRE_75 = 32'h00000000;
	wire [31:0] _regs_WIRE_76 = 32'h00000000;
	wire [31:0] _regs_WIRE_77 = 32'h00000000;
	wire [31:0] _regs_WIRE_78 = 32'h00000000;
	wire [31:0] _regs_WIRE_79 = 32'h00000000;
	wire [31:0] _regs_WIRE_80 = 32'h00000000;
	wire [31:0] _regs_WIRE_81 = 32'h00000000;
	wire [31:0] _regs_WIRE_82 = 32'h00000000;
	wire [31:0] _regs_WIRE_83 = 32'h00000000;
	wire [31:0] _regs_WIRE_84 = 32'h00000000;
	wire [31:0] _regs_WIRE_85 = 32'h00000000;
	wire [31:0] _regs_WIRE_86 = 32'h00000000;
	wire [31:0] _regs_WIRE_87 = 32'h00000000;
	wire [31:0] _regs_WIRE_88 = 32'h00000000;
	wire [31:0] _regs_WIRE_89 = 32'h00000000;
	wire [31:0] _regs_WIRE_90 = 32'h00000000;
	wire [31:0] _regs_WIRE_91 = 32'h00000000;
	wire [31:0] _regs_WIRE_92 = 32'h00000000;
	wire [31:0] _regs_WIRE_93 = 32'h00000000;
	wire [31:0] _regs_WIRE_94 = 32'h00000000;
	wire [31:0] _regs_WIRE_95 = 32'h00000000;
	wire [31:0] _regs_WIRE_96 = 32'h00000000;
	wire [31:0] _regs_WIRE_97 = 32'h00000000;
	wire [31:0] _regs_WIRE_98 = 32'h00000000;
	wire [31:0] _regs_WIRE_99 = 32'h00000000;
	wire [31:0] _regs_WIRE_100 = 32'h00000000;
	wire [31:0] _regs_WIRE_101 = 32'h00000000;
	wire [31:0] _regs_WIRE_102 = 32'h00000000;
	wire [31:0] _regs_WIRE_103 = 32'h00000000;
	wire [31:0] _regs_WIRE_104 = 32'h00000000;
	wire [31:0] _regs_WIRE_105 = 32'h00000000;
	wire [31:0] _regs_WIRE_106 = 32'h00000000;
	wire [31:0] _regs_WIRE_107 = 32'h00000000;
	wire [31:0] _regs_WIRE_108 = 32'h00000000;
	wire [31:0] _regs_WIRE_109 = 32'h00000000;
	wire [31:0] _regs_WIRE_110 = 32'h00000000;
	wire [31:0] _regs_WIRE_111 = 32'h00000000;
	wire [31:0] _regs_WIRE_112 = 32'h00000000;
	wire [31:0] _regs_WIRE_113 = 32'h00000000;
	wire [31:0] _regs_WIRE_114 = 32'h00000000;
	wire [31:0] _regs_WIRE_115 = 32'h00000000;
	wire [31:0] _regs_WIRE_116 = 32'h00000000;
	wire [31:0] _regs_WIRE_117 = 32'h00000000;
	wire [31:0] _regs_WIRE_118 = 32'h00000000;
	wire [31:0] _regs_WIRE_119 = 32'h00000000;
	wire [31:0] _regs_WIRE_120 = 32'h00000000;
	wire [31:0] _regs_WIRE_121 = 32'h00000000;
	wire [31:0] _regs_WIRE_122 = 32'h00000000;
	wire [31:0] _regs_WIRE_123 = 32'h00000000;
	wire [31:0] _regs_WIRE_124 = 32'h00000000;
	wire [31:0] _regs_WIRE_125 = 32'h00000000;
	wire [31:0] _regs_WIRE_126 = 32'h00000000;
	wire [31:0] _regs_WIRE_127 = 32'h00000000;
	reg [31:0] regs_0;
	reg [31:0] regs_1;
	reg [31:0] regs_2;
	reg [31:0] regs_3;
	reg [31:0] regs_4;
	reg [31:0] regs_5;
	reg [31:0] regs_6;
	reg [31:0] regs_7;
	reg [31:0] regs_8;
	reg [31:0] regs_9;
	reg [31:0] regs_10;
	reg [31:0] regs_11;
	reg [31:0] regs_12;
	reg [31:0] regs_13;
	reg [31:0] regs_14;
	reg [31:0] regs_15;
	reg [31:0] regs_16;
	reg [31:0] regs_17;
	reg [31:0] regs_18;
	reg [31:0] regs_19;
	reg [31:0] regs_20;
	reg [31:0] regs_21;
	reg [31:0] regs_22;
	reg [31:0] regs_23;
	reg [31:0] regs_24;
	reg [31:0] regs_25;
	reg [31:0] regs_26;
	reg [31:0] regs_27;
	reg [31:0] regs_28;
	reg [31:0] regs_29;
	reg [31:0] regs_30;
	reg [31:0] regs_31;
	reg [31:0] regs_32;
	reg [31:0] regs_33;
	reg [31:0] regs_34;
	reg [31:0] regs_35;
	reg [31:0] regs_36;
	reg [31:0] regs_37;
	reg [31:0] regs_38;
	reg [31:0] regs_39;
	reg [31:0] regs_40;
	reg [31:0] regs_41;
	reg [31:0] regs_42;
	reg [31:0] regs_43;
	reg [31:0] regs_44;
	reg [31:0] regs_45;
	reg [31:0] regs_46;
	reg [31:0] regs_47;
	reg [31:0] regs_48;
	reg [31:0] regs_49;
	reg [31:0] regs_50;
	reg [31:0] regs_51;
	reg [31:0] regs_52;
	reg [31:0] regs_53;
	reg [31:0] regs_54;
	reg [31:0] regs_55;
	reg [31:0] regs_56;
	reg [31:0] regs_57;
	reg [31:0] regs_58;
	reg [31:0] regs_59;
	reg [31:0] regs_60;
	reg [31:0] regs_61;
	reg [31:0] regs_62;
	reg [31:0] regs_63;
	reg [31:0] regs_64;
	reg [31:0] regs_65;
	reg [31:0] regs_66;
	reg [31:0] regs_67;
	reg [31:0] regs_68;
	reg [31:0] regs_69;
	reg [31:0] regs_70;
	reg [31:0] regs_71;
	reg [31:0] regs_72;
	reg [31:0] regs_73;
	reg [31:0] regs_74;
	reg [31:0] regs_75;
	reg [31:0] regs_76;
	reg [31:0] regs_77;
	reg [31:0] regs_78;
	reg [31:0] regs_79;
	reg [31:0] regs_80;
	reg [31:0] regs_81;
	reg [31:0] regs_82;
	reg [31:0] regs_83;
	reg [31:0] regs_84;
	reg [31:0] regs_85;
	reg [31:0] regs_86;
	reg [31:0] regs_87;
	reg [31:0] regs_88;
	reg [31:0] regs_89;
	reg [31:0] regs_90;
	reg [31:0] regs_91;
	reg [31:0] regs_92;
	reg [31:0] regs_93;
	reg [31:0] regs_94;
	reg [31:0] regs_95;
	reg [31:0] regs_96;
	reg [31:0] regs_97;
	reg [31:0] regs_98;
	reg [31:0] regs_99;
	reg [31:0] regs_100;
	reg [31:0] regs_101;
	reg [31:0] regs_102;
	reg [31:0] regs_103;
	reg [31:0] regs_104;
	reg [31:0] regs_105;
	reg [31:0] regs_106;
	reg [31:0] regs_107;
	reg [31:0] regs_108;
	reg [31:0] regs_109;
	reg [31:0] regs_110;
	reg [31:0] regs_111;
	reg [31:0] regs_112;
	reg [31:0] regs_113;
	reg [31:0] regs_114;
	reg [31:0] regs_115;
	reg [31:0] regs_116;
	reg [31:0] regs_117;
	reg [31:0] regs_118;
	reg [31:0] regs_119;
	reg [31:0] regs_120;
	reg [31:0] regs_121;
	reg [31:0] regs_122;
	reg [31:0] regs_123;
	reg [31:0] regs_124;
	reg [31:0] regs_125;
	reg [31:0] regs_126;
	reg [31:0] regs_127;
	wire [6:0] effectiveSrc1 = {io_threadID_0, io_src1_0};
	wire [6:0] effectiveSrc2 = {io_threadID_0, io_src2_0};
	wire [6:0] effectiveDst1 = {io_threadID_0, io_dst1_0};
	wire [4095:0] _GEN = {regs_127, regs_126, regs_125, regs_124, regs_123, regs_122, regs_121, regs_120, regs_119, regs_118, regs_117, regs_116, regs_115, regs_114, regs_113, regs_112, regs_111, regs_110, regs_109, regs_108, regs_107, regs_106, regs_105, regs_104, regs_103, regs_102, regs_101, regs_100, regs_99, regs_98, regs_97, regs_96, regs_95, regs_94, regs_93, regs_92, regs_91, regs_90, regs_89, regs_88, regs_87, regs_86, regs_85, regs_84, regs_83, regs_82, regs_81, regs_80, regs_79, regs_78, regs_77, regs_76, regs_75, regs_74, regs_73, regs_72, regs_71, regs_70, regs_69, regs_68, regs_67, regs_66, regs_65, regs_64, regs_63, regs_62, regs_61, regs_60, regs_59, regs_58, regs_57, regs_56, regs_55, regs_54, regs_53, regs_52, regs_51, regs_50, regs_49, regs_48, regs_47, regs_46, regs_45, regs_44, regs_43, regs_42, regs_41, regs_40, regs_39, regs_38, regs_37, regs_36, regs_35, regs_34, regs_33, regs_32, regs_31, regs_30, regs_29, regs_28, regs_27, regs_26, regs_25, regs_24, regs_23, regs_22, regs_21, regs_20, regs_19, regs_18, regs_17, regs_16, regs_15, regs_14, regs_13, regs_12, regs_11, regs_10, regs_9, regs_8, regs_7, regs_6, regs_5, regs_4, regs_3, regs_2, regs_1, regs_0};
	wire [31:0] io_src1data_0 = _GEN[effectiveSrc1 * 32+:32];
	wire [31:0] io_src2data_0 = _GEN[effectiveSrc2 * 32+:32];
	always @(posedge clock)
		if (reset) begin
			regs_0 <= 32'h00000000;
			regs_1 <= 32'h00000000;
			regs_2 <= 32'h00000000;
			regs_3 <= 32'h00000000;
			regs_4 <= 32'h00000000;
			regs_5 <= 32'h00000000;
			regs_6 <= 32'h00000000;
			regs_7 <= 32'h00000000;
			regs_8 <= 32'h00000000;
			regs_9 <= 32'h00000000;
			regs_10 <= 32'h00000000;
			regs_11 <= 32'h00000000;
			regs_12 <= 32'h00000000;
			regs_13 <= 32'h00000000;
			regs_14 <= 32'h00000000;
			regs_15 <= 32'h00000000;
			regs_16 <= 32'h00000000;
			regs_17 <= 32'h00000000;
			regs_18 <= 32'h00000000;
			regs_19 <= 32'h00000000;
			regs_20 <= 32'h00000000;
			regs_21 <= 32'h00000000;
			regs_22 <= 32'h00000000;
			regs_23 <= 32'h00000000;
			regs_24 <= 32'h00000000;
			regs_25 <= 32'h00000000;
			regs_26 <= 32'h00000000;
			regs_27 <= 32'h00000000;
			regs_28 <= 32'h00000000;
			regs_29 <= 32'h00000000;
			regs_30 <= 32'h00000000;
			regs_31 <= 32'h00000000;
			regs_32 <= 32'h00000000;
			regs_33 <= 32'h00000000;
			regs_34 <= 32'h00000000;
			regs_35 <= 32'h00000000;
			regs_36 <= 32'h00000000;
			regs_37 <= 32'h00000000;
			regs_38 <= 32'h00000000;
			regs_39 <= 32'h00000000;
			regs_40 <= 32'h00000000;
			regs_41 <= 32'h00000000;
			regs_42 <= 32'h00000000;
			regs_43 <= 32'h00000000;
			regs_44 <= 32'h00000000;
			regs_45 <= 32'h00000000;
			regs_46 <= 32'h00000000;
			regs_47 <= 32'h00000000;
			regs_48 <= 32'h00000000;
			regs_49 <= 32'h00000000;
			regs_50 <= 32'h00000000;
			regs_51 <= 32'h00000000;
			regs_52 <= 32'h00000000;
			regs_53 <= 32'h00000000;
			regs_54 <= 32'h00000000;
			regs_55 <= 32'h00000000;
			regs_56 <= 32'h00000000;
			regs_57 <= 32'h00000000;
			regs_58 <= 32'h00000000;
			regs_59 <= 32'h00000000;
			regs_60 <= 32'h00000000;
			regs_61 <= 32'h00000000;
			regs_62 <= 32'h00000000;
			regs_63 <= 32'h00000000;
			regs_64 <= 32'h00000000;
			regs_65 <= 32'h00000000;
			regs_66 <= 32'h00000000;
			regs_67 <= 32'h00000000;
			regs_68 <= 32'h00000000;
			regs_69 <= 32'h00000000;
			regs_70 <= 32'h00000000;
			regs_71 <= 32'h00000000;
			regs_72 <= 32'h00000000;
			regs_73 <= 32'h00000000;
			regs_74 <= 32'h00000000;
			regs_75 <= 32'h00000000;
			regs_76 <= 32'h00000000;
			regs_77 <= 32'h00000000;
			regs_78 <= 32'h00000000;
			regs_79 <= 32'h00000000;
			regs_80 <= 32'h00000000;
			regs_81 <= 32'h00000000;
			regs_82 <= 32'h00000000;
			regs_83 <= 32'h00000000;
			regs_84 <= 32'h00000000;
			regs_85 <= 32'h00000000;
			regs_86 <= 32'h00000000;
			regs_87 <= 32'h00000000;
			regs_88 <= 32'h00000000;
			regs_89 <= 32'h00000000;
			regs_90 <= 32'h00000000;
			regs_91 <= 32'h00000000;
			regs_92 <= 32'h00000000;
			regs_93 <= 32'h00000000;
			regs_94 <= 32'h00000000;
			regs_95 <= 32'h00000000;
			regs_96 <= 32'h00000000;
			regs_97 <= 32'h00000000;
			regs_98 <= 32'h00000000;
			regs_99 <= 32'h00000000;
			regs_100 <= 32'h00000000;
			regs_101 <= 32'h00000000;
			regs_102 <= 32'h00000000;
			regs_103 <= 32'h00000000;
			regs_104 <= 32'h00000000;
			regs_105 <= 32'h00000000;
			regs_106 <= 32'h00000000;
			regs_107 <= 32'h00000000;
			regs_108 <= 32'h00000000;
			regs_109 <= 32'h00000000;
			regs_110 <= 32'h00000000;
			regs_111 <= 32'h00000000;
			regs_112 <= 32'h00000000;
			regs_113 <= 32'h00000000;
			regs_114 <= 32'h00000000;
			regs_115 <= 32'h00000000;
			regs_116 <= 32'h00000000;
			regs_117 <= 32'h00000000;
			regs_118 <= 32'h00000000;
			regs_119 <= 32'h00000000;
			regs_120 <= 32'h00000000;
			regs_121 <= 32'h00000000;
			regs_122 <= 32'h00000000;
			regs_123 <= 32'h00000000;
			regs_124 <= 32'h00000000;
			regs_125 <= 32'h00000000;
			regs_126 <= 32'h00000000;
			regs_127 <= 32'h00000000;
		end
		else begin
			if (io_wen_0 & (effectiveDst1 == 7'h00))
				regs_0 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h01))
				regs_1 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h02))
				regs_2 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h03))
				regs_3 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h04))
				regs_4 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h05))
				regs_5 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h06))
				regs_6 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h07))
				regs_7 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h08))
				regs_8 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h09))
				regs_9 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h0a))
				regs_10 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h0b))
				regs_11 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h0c))
				regs_12 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h0d))
				regs_13 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h0e))
				regs_14 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h0f))
				regs_15 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h10))
				regs_16 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h11))
				regs_17 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h12))
				regs_18 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h13))
				regs_19 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h14))
				regs_20 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h15))
				regs_21 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h16))
				regs_22 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h17))
				regs_23 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h18))
				regs_24 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h19))
				regs_25 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h1a))
				regs_26 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h1b))
				regs_27 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h1c))
				regs_28 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h1d))
				regs_29 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h1e))
				regs_30 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h1f))
				regs_31 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h20))
				regs_32 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h21))
				regs_33 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h22))
				regs_34 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h23))
				regs_35 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h24))
				regs_36 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h25))
				regs_37 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h26))
				regs_38 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h27))
				regs_39 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h28))
				regs_40 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h29))
				regs_41 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h2a))
				regs_42 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h2b))
				regs_43 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h2c))
				regs_44 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h2d))
				regs_45 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h2e))
				regs_46 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h2f))
				regs_47 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h30))
				regs_48 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h31))
				regs_49 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h32))
				regs_50 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h33))
				regs_51 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h34))
				regs_52 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h35))
				regs_53 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h36))
				regs_54 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h37))
				regs_55 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h38))
				regs_56 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h39))
				regs_57 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h3a))
				regs_58 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h3b))
				regs_59 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h3c))
				regs_60 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h3d))
				regs_61 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h3e))
				regs_62 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h3f))
				regs_63 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h40))
				regs_64 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h41))
				regs_65 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h42))
				regs_66 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h43))
				regs_67 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h44))
				regs_68 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h45))
				regs_69 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h46))
				regs_70 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h47))
				regs_71 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h48))
				regs_72 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h49))
				regs_73 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h4a))
				regs_74 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h4b))
				regs_75 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h4c))
				regs_76 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h4d))
				regs_77 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h4e))
				regs_78 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h4f))
				regs_79 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h50))
				regs_80 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h51))
				regs_81 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h52))
				regs_82 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h53))
				regs_83 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h54))
				regs_84 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h55))
				regs_85 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h56))
				regs_86 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h57))
				regs_87 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h58))
				regs_88 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h59))
				regs_89 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h5a))
				regs_90 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h5b))
				regs_91 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h5c))
				regs_92 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h5d))
				regs_93 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h5e))
				regs_94 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h5f))
				regs_95 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h60))
				regs_96 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h61))
				regs_97 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h62))
				regs_98 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h63))
				regs_99 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h64))
				regs_100 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h65))
				regs_101 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h66))
				regs_102 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h67))
				regs_103 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h68))
				regs_104 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h69))
				regs_105 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h6a))
				regs_106 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h6b))
				regs_107 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h6c))
				regs_108 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h6d))
				regs_109 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h6e))
				regs_110 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h6f))
				regs_111 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h70))
				regs_112 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h71))
				regs_113 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h72))
				regs_114 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h73))
				regs_115 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h74))
				regs_116 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h75))
				regs_117 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h76))
				regs_118 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h77))
				regs_119 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h78))
				regs_120 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h79))
				regs_121 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h7a))
				regs_122 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h7b))
				regs_123 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h7c))
				regs_124 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h7d))
				regs_125 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h7e))
				regs_126 <= io_dst1data_0;
			if (io_wen_0 & (&effectiveDst1))
				regs_127 <= io_dst1data_0;
		end
	initial begin : sv2v_autoblock_1
		reg [31:0] _RANDOM [0:127];
	end
	assign io_src1data = io_src1data_0;
	assign io_src2data = io_src2data_0;
endmodule
