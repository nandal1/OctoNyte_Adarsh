module RISCVAdderSubtractor32 (
	clock,
	reset,
	io_a,
	io_b,
	io_opcode,
	io_carryIn,
	io_result,
	io_carryOut,
	io_overflowFlag,
	io_zeroFlag,
	io_negativeFlag
);
	input clock;
	input reset;
	input [31:0] io_a;
	input [31:0] io_b;
	input [3:0] io_opcode;
	input io_carryIn;
	output wire [31:0] io_result;
	output wire io_carryOut;
	output wire io_overflowFlag;
	output wire io_zeroFlag;
	output wire io_negativeFlag;
	wire [31:0] io_a_0 = io_a;
	wire [31:0] io_b_0 = io_b;
	wire [3:0] io_opcode_0 = io_opcode;
	wire io_carryIn_0 = io_carryIn;
	wire [5:0] _width_T_3 = 6'h20;
	wire [31:0] _mask_T_3 = 32'hffffffff;
	wire _io_carryOut_T_6;
	wire isOverflow;
	wire isZero;
	wire isNegative;
	wire _isSub_T = io_opcode_0[3];
	wire isSub = _isSub_T;
	wire isSigned = io_opcode_0[2];
	wire [1:0] operandSize = io_opcode_0[1:0];
	wire _GEN = operandSize == 2'h0;
	wire _width_T;
	assign _width_T = _GEN;
	wire _mask_T;
	assign _mask_T = _GEN;
	wire _GEN_0 = operandSize == 2'h1;
	wire _width_T_1;
	assign _width_T_1 = _GEN_0;
	wire _mask_T_1;
	assign _mask_T_1 = _GEN_0;
	wire _GEN_1 = operandSize == 2'h2;
	wire _width_T_2;
	assign _width_T_2 = _GEN_1;
	wire _mask_T_2;
	assign _mask_T_2 = _GEN_1;
	wire [5:0] _width_T_4 = (_width_T_1 ? 6'h10 : 6'h20);
	wire [5:0] width = (_width_T ? 6'h08 : _width_T_4);
	wire [31:0] _mask_T_4 = (_mask_T_1 ? 32'h0000ffff : 32'hffffffff);
	wire [31:0] mask = (_mask_T ? 32'h000000ff : _mask_T_4);
	wire [31:0] aEffective = io_a_0 & mask;
	wire [31:0] _fullArithmeticResult_T = aEffective;
	wire [31:0] bEffective = io_b_0 & mask;
	wire [31:0] _bAdjusted_T = ~bEffective;
	wire [32:0] _bAdjusted_T_1 = {1'h0, _bAdjusted_T} + 33'h000000001;
	wire [31:0] _bAdjusted_T_2 = _bAdjusted_T_1[31:0];
	wire [31:0] bAdjusted = (isSub ? _bAdjusted_T_2 : bEffective);
	wire [31:0] _fullArithmeticResult_T_1 = bAdjusted;
	wire [32:0] _fullArithmeticResult_T_2 = {_fullArithmeticResult_T[31], _fullArithmeticResult_T} + {_fullArithmeticResult_T_1[31], _fullArithmeticResult_T_1};
	wire [32:0] _fullArithmeticResult_T_3 = _fullArithmeticResult_T_2;
	wire [32:0] _fullArithmeticResult_T_4 = {1'h0, aEffective} + {1'h0, bAdjusted};
	wire [32:0] fullArithmeticResult = (isSigned ? _fullArithmeticResult_T_3 : _fullArithmeticResult_T_4);
	wire [32:0] truncatedResult = {1'h0, fullArithmeticResult[31:0] & mask};
	wire [31:0] io_result_0 = truncatedResult[31:0];
	wire _GEN_2 = width == 6'h08;
	wire _isCarry_T;
	assign _isCarry_T = _GEN_2;
	wire _aSign_T;
	assign _aSign_T = _GEN_2;
	wire _bSign_T;
	assign _bSign_T = _GEN_2;
	wire _sumSign_T;
	assign _sumSign_T = _GEN_2;
	wire _isCarry_T_1 = fullArithmeticResult[8];
	wire _GEN_3 = width == 6'h10;
	wire _isCarry_T_2;
	assign _isCarry_T_2 = _GEN_3;
	wire _aSign_T_2;
	assign _aSign_T_2 = _GEN_3;
	wire _bSign_T_2;
	assign _bSign_T_2 = _GEN_3;
	wire _sumSign_T_2;
	assign _sumSign_T_2 = _GEN_3;
	wire _isCarry_T_3 = fullArithmeticResult[16];
	wire _GEN_4 = width == 6'h20;
	wire _isCarry_T_4;
	assign _isCarry_T_4 = _GEN_4;
	wire _aSign_T_4;
	assign _aSign_T_4 = _GEN_4;
	wire _bSign_T_4;
	assign _bSign_T_4 = _GEN_4;
	wire _sumSign_T_4;
	assign _sumSign_T_4 = _GEN_4;
	wire _isCarry_T_5 = fullArithmeticResult[32];
	wire _isCarry_T_6 = _isCarry_T_4 & _isCarry_T_5;
	wire _isCarry_T_7 = (_isCarry_T_2 ? _isCarry_T_3 : _isCarry_T_6);
	wire isCarry = (_isCarry_T ? _isCarry_T_1 : _isCarry_T_7);
	wire _isBorrow_T = ~isSigned;
	wire _isBorrow_T_1 = isSub & _isBorrow_T;
	wire _isBorrow_T_2 = aEffective < bEffective;
	wire isBorrow = _isBorrow_T_1 & _isBorrow_T_2;
	wire _io_carryOut_T = ~isSigned;
	wire _io_carryOut_T_1 = ~isSub;
	wire _io_carryOut_T_2 = _io_carryOut_T & _io_carryOut_T_1;
	wire _io_carryOut_T_3 = ~isSigned;
	wire _io_carryOut_T_4 = _io_carryOut_T_3 & isSub;
	wire _io_carryOut_T_5 = _io_carryOut_T_4 & isBorrow;
	assign _io_carryOut_T_6 = (_io_carryOut_T_2 ? isCarry : _io_carryOut_T_5);
	wire io_carryOut_0 = _io_carryOut_T_6;
	wire _aSign_T_8;
	wire _bSign_T_8;
	wire _sumSign_T_8;
	wire _aSign_T_1 = aEffective[7];
	wire _aSign_T_3 = aEffective[15];
	wire _aSign_T_5 = aEffective[31];
	wire _aSign_T_6 = _aSign_T_4 & _aSign_T_5;
	wire _aSign_T_7 = (_aSign_T_2 ? _aSign_T_3 : _aSign_T_6);
	assign _aSign_T_8 = (_aSign_T ? _aSign_T_1 : _aSign_T_7);
	wire aSign = _aSign_T_8;
	wire _bSign_T_1 = bAdjusted[7];
	wire _bSign_T_3 = bAdjusted[15];
	wire _bSign_T_5 = bAdjusted[31];
	wire _bSign_T_6 = _bSign_T_4 & _bSign_T_5;
	wire _bSign_T_7 = (_bSign_T_2 ? _bSign_T_3 : _bSign_T_6);
	assign _bSign_T_8 = (_bSign_T ? _bSign_T_1 : _bSign_T_7);
	wire bSign = _bSign_T_8;
	wire _sumSign_T_1 = fullArithmeticResult[7];
	wire _sumSign_T_3 = fullArithmeticResult[15];
	wire _sumSign_T_5 = fullArithmeticResult[31];
	wire _sumSign_T_6 = _sumSign_T_4 & _sumSign_T_5;
	wire _sumSign_T_7 = (_sumSign_T_2 ? _sumSign_T_3 : _sumSign_T_6);
	assign _sumSign_T_8 = (_sumSign_T ? _sumSign_T_1 : _sumSign_T_7);
	wire sumSign = _sumSign_T_8;
	wire _isOverflow_T = aSign == bSign;
	wire _isOverflow_T_1 = aSign != sumSign;
	assign isOverflow = _isOverflow_T & _isOverflow_T_1;
	wire io_overflowFlag_0 = isOverflow;
	wire _isZero_T = |truncatedResult;
	assign isZero = ~_isZero_T;
	wire io_zeroFlag_0 = isZero;
	assign isNegative = isSigned & sumSign;
	wire io_negativeFlag_0 = isNegative;
	assign io_result = io_result_0;
	assign io_carryOut = io_carryOut_0;
	assign io_overflowFlag = io_overflowFlag_0;
	assign io_zeroFlag = io_zeroFlag_0;
	assign io_negativeFlag = io_negativeFlag_0;
endmodule
