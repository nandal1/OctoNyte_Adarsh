module RegFileMT2R1WVec (
	clock,
	reset,
	io_threadID,
	io_src1,
	io_src2,
	io_dst1,
	io_wen,
	io_dst1data,
	io_src1data,
	io_src2data
);
	input clock;
	input reset;
	input [1:0] io_threadID;
	input [4:0] io_src1;
	input [4:0] io_src2;
	input [4:0] io_dst1;
	input io_wen;
	input [31:0] io_dst1data;
	output wire [31:0] io_src1data;
	output wire [31:0] io_src2data;
	wire [1:0] io_threadID_0 = io_threadID;
	wire [4:0] io_src1_0 = io_src1;
	wire [4:0] io_src2_0 = io_src2;
	wire [4:0] io_dst1_0 = io_dst1;
	wire io_wen_0 = io_wen;
	wire [31:0] io_dst1data_0 = io_dst1data;
	wire [31:0] _regs_WIRE_0 = 32'h00000000;
	wire [31:0] _regs_WIRE_1 = 32'h00000000;
	wire [31:0] _regs_WIRE_2 = 32'h00000000;
	wire [31:0] _regs_WIRE_3 = 32'h00000000;
	wire [31:0] _regs_WIRE_4 = 32'h00000000;
	wire [31:0] _regs_WIRE_5 = 32'h00000000;
	wire [31:0] _regs_WIRE_6 = 32'h00000000;
	wire [31:0] _regs_WIRE_7 = 32'h00000000;
	wire [31:0] _regs_WIRE_8 = 32'h00000000;
	wire [31:0] _regs_WIRE_9 = 32'h00000000;
	wire [31:0] _regs_WIRE_10 = 32'h00000000;
	wire [31:0] _regs_WIRE_11 = 32'h00000000;
	wire [31:0] _regs_WIRE_12 = 32'h00000000;
	wire [31:0] _regs_WIRE_13 = 32'h00000000;
	wire [31:0] _regs_WIRE_14 = 32'h00000000;
	wire [31:0] _regs_WIRE_15 = 32'h00000000;
	wire [31:0] _regs_WIRE_16 = 32'h00000000;
	wire [31:0] _regs_WIRE_17 = 32'h00000000;
	wire [31:0] _regs_WIRE_18 = 32'h00000000;
	wire [31:0] _regs_WIRE_19 = 32'h00000000;
	wire [31:0] _regs_WIRE_20 = 32'h00000000;
	wire [31:0] _regs_WIRE_21 = 32'h00000000;
	wire [31:0] _regs_WIRE_22 = 32'h00000000;
	wire [31:0] _regs_WIRE_23 = 32'h00000000;
	wire [31:0] _regs_WIRE_24 = 32'h00000000;
	wire [31:0] _regs_WIRE_25 = 32'h00000000;
	wire [31:0] _regs_WIRE_26 = 32'h00000000;
	wire [31:0] _regs_WIRE_27 = 32'h00000000;
	wire [31:0] _regs_WIRE_28 = 32'h00000000;
	wire [31:0] _regs_WIRE_29 = 32'h00000000;
	wire [31:0] _regs_WIRE_30 = 32'h00000000;
	wire [31:0] _regs_WIRE_31 = 32'h00000000;
	wire [31:0] _regs_WIRE_32 = 32'h00000000;
	wire [31:0] _regs_WIRE_33 = 32'h00000000;
	wire [31:0] _regs_WIRE_34 = 32'h00000000;
	wire [31:0] _regs_WIRE_35 = 32'h00000000;
	wire [31:0] _regs_WIRE_36 = 32'h00000000;
	wire [31:0] _regs_WIRE_37 = 32'h00000000;
	wire [31:0] _regs_WIRE_38 = 32'h00000000;
	wire [31:0] _regs_WIRE_39 = 32'h00000000;
	wire [31:0] _regs_WIRE_40 = 32'h00000000;
	wire [31:0] _regs_WIRE_41 = 32'h00000000;
	wire [31:0] _regs_WIRE_42 = 32'h00000000;
	wire [31:0] _regs_WIRE_43 = 32'h00000000;
	wire [31:0] _regs_WIRE_44 = 32'h00000000;
	wire [31:0] _regs_WIRE_45 = 32'h00000000;
	wire [31:0] _regs_WIRE_46 = 32'h00000000;
	wire [31:0] _regs_WIRE_47 = 32'h00000000;
	wire [31:0] _regs_WIRE_48 = 32'h00000000;
	wire [31:0] _regs_WIRE_49 = 32'h00000000;
	wire [31:0] _regs_WIRE_50 = 32'h00000000;
	wire [31:0] _regs_WIRE_51 = 32'h00000000;
	wire [31:0] _regs_WIRE_52 = 32'h00000000;
	wire [31:0] _regs_WIRE_53 = 32'h00000000;
	wire [31:0] _regs_WIRE_54 = 32'h00000000;
	wire [31:0] _regs_WIRE_55 = 32'h00000000;
	wire [31:0] _regs_WIRE_56 = 32'h00000000;
	wire [31:0] _regs_WIRE_57 = 32'h00000000;
	wire [31:0] _regs_WIRE_58 = 32'h00000000;
	wire [31:0] _regs_WIRE_59 = 32'h00000000;
	wire [31:0] _regs_WIRE_60 = 32'h00000000;
	wire [31:0] _regs_WIRE_61 = 32'h00000000;
	wire [31:0] _regs_WIRE_62 = 32'h00000000;
	wire [31:0] _regs_WIRE_63 = 32'h00000000;
	wire [31:0] _regs_WIRE_64 = 32'h00000000;
	wire [31:0] _regs_WIRE_65 = 32'h00000000;
	wire [31:0] _regs_WIRE_66 = 32'h00000000;
	wire [31:0] _regs_WIRE_67 = 32'h00000000;
	wire [31:0] _regs_WIRE_68 = 32'h00000000;
	wire [31:0] _regs_WIRE_69 = 32'h00000000;
	wire [31:0] _regs_WIRE_70 = 32'h00000000;
	wire [31:0] _regs_WIRE_71 = 32'h00000000;
	wire [31:0] _regs_WIRE_72 = 32'h00000000;
	wire [31:0] _regs_WIRE_73 = 32'h00000000;
	wire [31:0] _regs_WIRE_74 = 32'h00000000;
	wire [31:0] _regs_WIRE_75 = 32'h00000000;
	wire [31:0] _regs_WIRE_76 = 32'h00000000;
	wire [31:0] _regs_WIRE_77 = 32'h00000000;
	wire [31:0] _regs_WIRE_78 = 32'h00000000;
	wire [31:0] _regs_WIRE_79 = 32'h00000000;
	wire [31:0] _regs_WIRE_80 = 32'h00000000;
	wire [31:0] _regs_WIRE_81 = 32'h00000000;
	wire [31:0] _regs_WIRE_82 = 32'h00000000;
	wire [31:0] _regs_WIRE_83 = 32'h00000000;
	wire [31:0] _regs_WIRE_84 = 32'h00000000;
	wire [31:0] _regs_WIRE_85 = 32'h00000000;
	wire [31:0] _regs_WIRE_86 = 32'h00000000;
	wire [31:0] _regs_WIRE_87 = 32'h00000000;
	wire [31:0] _regs_WIRE_88 = 32'h00000000;
	wire [31:0] _regs_WIRE_89 = 32'h00000000;
	wire [31:0] _regs_WIRE_90 = 32'h00000000;
	wire [31:0] _regs_WIRE_91 = 32'h00000000;
	wire [31:0] _regs_WIRE_92 = 32'h00000000;
	wire [31:0] _regs_WIRE_93 = 32'h00000000;
	wire [31:0] _regs_WIRE_94 = 32'h00000000;
	wire [31:0] _regs_WIRE_95 = 32'h00000000;
	wire [31:0] _regs_WIRE_96 = 32'h00000000;
	wire [31:0] _regs_WIRE_97 = 32'h00000000;
	wire [31:0] _regs_WIRE_98 = 32'h00000000;
	wire [31:0] _regs_WIRE_99 = 32'h00000000;
	wire [31:0] _regs_WIRE_100 = 32'h00000000;
	wire [31:0] _regs_WIRE_101 = 32'h00000000;
	wire [31:0] _regs_WIRE_102 = 32'h00000000;
	wire [31:0] _regs_WIRE_103 = 32'h00000000;
	wire [31:0] _regs_WIRE_104 = 32'h00000000;
	wire [31:0] _regs_WIRE_105 = 32'h00000000;
	wire [31:0] _regs_WIRE_106 = 32'h00000000;
	wire [31:0] _regs_WIRE_107 = 32'h00000000;
	wire [31:0] _regs_WIRE_108 = 32'h00000000;
	wire [31:0] _regs_WIRE_109 = 32'h00000000;
	wire [31:0] _regs_WIRE_110 = 32'h00000000;
	wire [31:0] _regs_WIRE_111 = 32'h00000000;
	wire [31:0] _regs_WIRE_112 = 32'h00000000;
	wire [31:0] _regs_WIRE_113 = 32'h00000000;
	wire [31:0] _regs_WIRE_114 = 32'h00000000;
	wire [31:0] _regs_WIRE_115 = 32'h00000000;
	wire [31:0] _regs_WIRE_116 = 32'h00000000;
	wire [31:0] _regs_WIRE_117 = 32'h00000000;
	wire [31:0] _regs_WIRE_118 = 32'h00000000;
	wire [31:0] _regs_WIRE_119 = 32'h00000000;
	wire [31:0] _regs_WIRE_120 = 32'h00000000;
	wire [31:0] _regs_WIRE_121 = 32'h00000000;
	wire [31:0] _regs_WIRE_122 = 32'h00000000;
	wire [31:0] _regs_WIRE_123 = 32'h00000000;
	wire [31:0] _regs_WIRE_124 = 32'h00000000;
	wire [31:0] _regs_WIRE_125 = 32'h00000000;
	wire [31:0] _regs_WIRE_126 = 32'h00000000;
	wire [31:0] _regs_WIRE_127 = 32'h00000000;
	reg [31:0] regs_0;
	reg [31:0] regs_1;
	reg [31:0] regs_2;
	reg [31:0] regs_3;
	reg [31:0] regs_4;
	reg [31:0] regs_5;
	reg [31:0] regs_6;
	reg [31:0] regs_7;
	reg [31:0] regs_8;
	reg [31:0] regs_9;
	reg [31:0] regs_10;
	reg [31:0] regs_11;
	reg [31:0] regs_12;
	reg [31:0] regs_13;
	reg [31:0] regs_14;
	reg [31:0] regs_15;
	reg [31:0] regs_16;
	reg [31:0] regs_17;
	reg [31:0] regs_18;
	reg [31:0] regs_19;
	reg [31:0] regs_20;
	reg [31:0] regs_21;
	reg [31:0] regs_22;
	reg [31:0] regs_23;
	reg [31:0] regs_24;
	reg [31:0] regs_25;
	reg [31:0] regs_26;
	reg [31:0] regs_27;
	reg [31:0] regs_28;
	reg [31:0] regs_29;
	reg [31:0] regs_30;
	reg [31:0] regs_31;
	reg [31:0] regs_32;
	reg [31:0] regs_33;
	reg [31:0] regs_34;
	reg [31:0] regs_35;
	reg [31:0] regs_36;
	reg [31:0] regs_37;
	reg [31:0] regs_38;
	reg [31:0] regs_39;
	reg [31:0] regs_40;
	reg [31:0] regs_41;
	reg [31:0] regs_42;
	reg [31:0] regs_43;
	reg [31:0] regs_44;
	reg [31:0] regs_45;
	reg [31:0] regs_46;
	reg [31:0] regs_47;
	reg [31:0] regs_48;
	reg [31:0] regs_49;
	reg [31:0] regs_50;
	reg [31:0] regs_51;
	reg [31:0] regs_52;
	reg [31:0] regs_53;
	reg [31:0] regs_54;
	reg [31:0] regs_55;
	reg [31:0] regs_56;
	reg [31:0] regs_57;
	reg [31:0] regs_58;
	reg [31:0] regs_59;
	reg [31:0] regs_60;
	reg [31:0] regs_61;
	reg [31:0] regs_62;
	reg [31:0] regs_63;
	reg [31:0] regs_64;
	reg [31:0] regs_65;
	reg [31:0] regs_66;
	reg [31:0] regs_67;
	reg [31:0] regs_68;
	reg [31:0] regs_69;
	reg [31:0] regs_70;
	reg [31:0] regs_71;
	reg [31:0] regs_72;
	reg [31:0] regs_73;
	reg [31:0] regs_74;
	reg [31:0] regs_75;
	reg [31:0] regs_76;
	reg [31:0] regs_77;
	reg [31:0] regs_78;
	reg [31:0] regs_79;
	reg [31:0] regs_80;
	reg [31:0] regs_81;
	reg [31:0] regs_82;
	reg [31:0] regs_83;
	reg [31:0] regs_84;
	reg [31:0] regs_85;
	reg [31:0] regs_86;
	reg [31:0] regs_87;
	reg [31:0] regs_88;
	reg [31:0] regs_89;
	reg [31:0] regs_90;
	reg [31:0] regs_91;
	reg [31:0] regs_92;
	reg [31:0] regs_93;
	reg [31:0] regs_94;
	reg [31:0] regs_95;
	reg [31:0] regs_96;
	reg [31:0] regs_97;
	reg [31:0] regs_98;
	reg [31:0] regs_99;
	reg [31:0] regs_100;
	reg [31:0] regs_101;
	reg [31:0] regs_102;
	reg [31:0] regs_103;
	reg [31:0] regs_104;
	reg [31:0] regs_105;
	reg [31:0] regs_106;
	reg [31:0] regs_107;
	reg [31:0] regs_108;
	reg [31:0] regs_109;
	reg [31:0] regs_110;
	reg [31:0] regs_111;
	reg [31:0] regs_112;
	reg [31:0] regs_113;
	reg [31:0] regs_114;
	reg [31:0] regs_115;
	reg [31:0] regs_116;
	reg [31:0] regs_117;
	reg [31:0] regs_118;
	reg [31:0] regs_119;
	reg [31:0] regs_120;
	reg [31:0] regs_121;
	reg [31:0] regs_122;
	reg [31:0] regs_123;
	reg [31:0] regs_124;
	reg [31:0] regs_125;
	reg [31:0] regs_126;
	reg [31:0] regs_127;
	wire [6:0] effectiveSrc1 = {io_threadID_0, io_src1_0};
	wire [6:0] effectiveSrc2 = {io_threadID_0, io_src2_0};
	wire [6:0] effectiveDst1 = {io_threadID_0, io_dst1_0};
	wire [4095:0] _GEN = {regs_127, regs_126, regs_125, regs_124, regs_123, regs_122, regs_121, regs_120, regs_119, regs_118, regs_117, regs_116, regs_115, regs_114, regs_113, regs_112, regs_111, regs_110, regs_109, regs_108, regs_107, regs_106, regs_105, regs_104, regs_103, regs_102, regs_101, regs_100, regs_99, regs_98, regs_97, regs_96, regs_95, regs_94, regs_93, regs_92, regs_91, regs_90, regs_89, regs_88, regs_87, regs_86, regs_85, regs_84, regs_83, regs_82, regs_81, regs_80, regs_79, regs_78, regs_77, regs_76, regs_75, regs_74, regs_73, regs_72, regs_71, regs_70, regs_69, regs_68, regs_67, regs_66, regs_65, regs_64, regs_63, regs_62, regs_61, regs_60, regs_59, regs_58, regs_57, regs_56, regs_55, regs_54, regs_53, regs_52, regs_51, regs_50, regs_49, regs_48, regs_47, regs_46, regs_45, regs_44, regs_43, regs_42, regs_41, regs_40, regs_39, regs_38, regs_37, regs_36, regs_35, regs_34, regs_33, regs_32, regs_31, regs_30, regs_29, regs_28, regs_27, regs_26, regs_25, regs_24, regs_23, regs_22, regs_21, regs_20, regs_19, regs_18, regs_17, regs_16, regs_15, regs_14, regs_13, regs_12, regs_11, regs_10, regs_9, regs_8, regs_7, regs_6, regs_5, regs_4, regs_3, regs_2, regs_1, regs_0};
	wire [31:0] io_src1data_0 = _GEN[effectiveSrc1 * 32+:32];
	wire [31:0] io_src2data_0 = _GEN[effectiveSrc2 * 32+:32];
	always @(posedge clock)
		if (reset) begin
			regs_0 <= 32'h00000000;
			regs_1 <= 32'h00000000;
			regs_2 <= 32'h00000000;
			regs_3 <= 32'h00000000;
			regs_4 <= 32'h00000000;
			regs_5 <= 32'h00000000;
			regs_6 <= 32'h00000000;
			regs_7 <= 32'h00000000;
			regs_8 <= 32'h00000000;
			regs_9 <= 32'h00000000;
			regs_10 <= 32'h00000000;
			regs_11 <= 32'h00000000;
			regs_12 <= 32'h00000000;
			regs_13 <= 32'h00000000;
			regs_14 <= 32'h00000000;
			regs_15 <= 32'h00000000;
			regs_16 <= 32'h00000000;
			regs_17 <= 32'h00000000;
			regs_18 <= 32'h00000000;
			regs_19 <= 32'h00000000;
			regs_20 <= 32'h00000000;
			regs_21 <= 32'h00000000;
			regs_22 <= 32'h00000000;
			regs_23 <= 32'h00000000;
			regs_24 <= 32'h00000000;
			regs_25 <= 32'h00000000;
			regs_26 <= 32'h00000000;
			regs_27 <= 32'h00000000;
			regs_28 <= 32'h00000000;
			regs_29 <= 32'h00000000;
			regs_30 <= 32'h00000000;
			regs_31 <= 32'h00000000;
			regs_32 <= 32'h00000000;
			regs_33 <= 32'h00000000;
			regs_34 <= 32'h00000000;
			regs_35 <= 32'h00000000;
			regs_36 <= 32'h00000000;
			regs_37 <= 32'h00000000;
			regs_38 <= 32'h00000000;
			regs_39 <= 32'h00000000;
			regs_40 <= 32'h00000000;
			regs_41 <= 32'h00000000;
			regs_42 <= 32'h00000000;
			regs_43 <= 32'h00000000;
			regs_44 <= 32'h00000000;
			regs_45 <= 32'h00000000;
			regs_46 <= 32'h00000000;
			regs_47 <= 32'h00000000;
			regs_48 <= 32'h00000000;
			regs_49 <= 32'h00000000;
			regs_50 <= 32'h00000000;
			regs_51 <= 32'h00000000;
			regs_52 <= 32'h00000000;
			regs_53 <= 32'h00000000;
			regs_54 <= 32'h00000000;
			regs_55 <= 32'h00000000;
			regs_56 <= 32'h00000000;
			regs_57 <= 32'h00000000;
			regs_58 <= 32'h00000000;
			regs_59 <= 32'h00000000;
			regs_60 <= 32'h00000000;
			regs_61 <= 32'h00000000;
			regs_62 <= 32'h00000000;
			regs_63 <= 32'h00000000;
			regs_64 <= 32'h00000000;
			regs_65 <= 32'h00000000;
			regs_66 <= 32'h00000000;
			regs_67 <= 32'h00000000;
			regs_68 <= 32'h00000000;
			regs_69 <= 32'h00000000;
			regs_70 <= 32'h00000000;
			regs_71 <= 32'h00000000;
			regs_72 <= 32'h00000000;
			regs_73 <= 32'h00000000;
			regs_74 <= 32'h00000000;
			regs_75 <= 32'h00000000;
			regs_76 <= 32'h00000000;
			regs_77 <= 32'h00000000;
			regs_78 <= 32'h00000000;
			regs_79 <= 32'h00000000;
			regs_80 <= 32'h00000000;
			regs_81 <= 32'h00000000;
			regs_82 <= 32'h00000000;
			regs_83 <= 32'h00000000;
			regs_84 <= 32'h00000000;
			regs_85 <= 32'h00000000;
			regs_86 <= 32'h00000000;
			regs_87 <= 32'h00000000;
			regs_88 <= 32'h00000000;
			regs_89 <= 32'h00000000;
			regs_90 <= 32'h00000000;
			regs_91 <= 32'h00000000;
			regs_92 <= 32'h00000000;
			regs_93 <= 32'h00000000;
			regs_94 <= 32'h00000000;
			regs_95 <= 32'h00000000;
			regs_96 <= 32'h00000000;
			regs_97 <= 32'h00000000;
			regs_98 <= 32'h00000000;
			regs_99 <= 32'h00000000;
			regs_100 <= 32'h00000000;
			regs_101 <= 32'h00000000;
			regs_102 <= 32'h00000000;
			regs_103 <= 32'h00000000;
			regs_104 <= 32'h00000000;
			regs_105 <= 32'h00000000;
			regs_106 <= 32'h00000000;
			regs_107 <= 32'h00000000;
			regs_108 <= 32'h00000000;
			regs_109 <= 32'h00000000;
			regs_110 <= 32'h00000000;
			regs_111 <= 32'h00000000;
			regs_112 <= 32'h00000000;
			regs_113 <= 32'h00000000;
			regs_114 <= 32'h00000000;
			regs_115 <= 32'h00000000;
			regs_116 <= 32'h00000000;
			regs_117 <= 32'h00000000;
			regs_118 <= 32'h00000000;
			regs_119 <= 32'h00000000;
			regs_120 <= 32'h00000000;
			regs_121 <= 32'h00000000;
			regs_122 <= 32'h00000000;
			regs_123 <= 32'h00000000;
			regs_124 <= 32'h00000000;
			regs_125 <= 32'h00000000;
			regs_126 <= 32'h00000000;
			regs_127 <= 32'h00000000;
		end
		else begin
			if (io_wen_0 & (effectiveDst1 == 7'h00))
				regs_0 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h01))
				regs_1 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h02))
				regs_2 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h03))
				regs_3 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h04))
				regs_4 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h05))
				regs_5 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h06))
				regs_6 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h07))
				regs_7 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h08))
				regs_8 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h09))
				regs_9 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h0a))
				regs_10 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h0b))
				regs_11 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h0c))
				regs_12 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h0d))
				regs_13 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h0e))
				regs_14 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h0f))
				regs_15 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h10))
				regs_16 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h11))
				regs_17 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h12))
				regs_18 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h13))
				regs_19 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h14))
				regs_20 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h15))
				regs_21 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h16))
				regs_22 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h17))
				regs_23 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h18))
				regs_24 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h19))
				regs_25 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h1a))
				regs_26 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h1b))
				regs_27 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h1c))
				regs_28 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h1d))
				regs_29 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h1e))
				regs_30 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h1f))
				regs_31 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h20))
				regs_32 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h21))
				regs_33 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h22))
				regs_34 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h23))
				regs_35 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h24))
				regs_36 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h25))
				regs_37 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h26))
				regs_38 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h27))
				regs_39 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h28))
				regs_40 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h29))
				regs_41 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h2a))
				regs_42 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h2b))
				regs_43 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h2c))
				regs_44 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h2d))
				regs_45 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h2e))
				regs_46 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h2f))
				regs_47 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h30))
				regs_48 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h31))
				regs_49 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h32))
				regs_50 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h33))
				regs_51 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h34))
				regs_52 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h35))
				regs_53 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h36))
				regs_54 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h37))
				regs_55 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h38))
				regs_56 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h39))
				regs_57 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h3a))
				regs_58 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h3b))
				regs_59 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h3c))
				regs_60 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h3d))
				regs_61 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h3e))
				regs_62 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h3f))
				regs_63 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h40))
				regs_64 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h41))
				regs_65 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h42))
				regs_66 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h43))
				regs_67 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h44))
				regs_68 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h45))
				regs_69 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h46))
				regs_70 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h47))
				regs_71 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h48))
				regs_72 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h49))
				regs_73 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h4a))
				regs_74 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h4b))
				regs_75 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h4c))
				regs_76 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h4d))
				regs_77 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h4e))
				regs_78 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h4f))
				regs_79 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h50))
				regs_80 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h51))
				regs_81 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h52))
				regs_82 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h53))
				regs_83 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h54))
				regs_84 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h55))
				regs_85 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h56))
				regs_86 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h57))
				regs_87 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h58))
				regs_88 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h59))
				regs_89 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h5a))
				regs_90 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h5b))
				regs_91 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h5c))
				regs_92 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h5d))
				regs_93 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h5e))
				regs_94 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h5f))
				regs_95 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h60))
				regs_96 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h61))
				regs_97 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h62))
				regs_98 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h63))
				regs_99 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h64))
				regs_100 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h65))
				regs_101 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h66))
				regs_102 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h67))
				regs_103 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h68))
				regs_104 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h69))
				regs_105 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h6a))
				regs_106 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h6b))
				regs_107 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h6c))
				regs_108 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h6d))
				regs_109 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h6e))
				regs_110 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h6f))
				regs_111 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h70))
				regs_112 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h71))
				regs_113 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h72))
				regs_114 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h73))
				regs_115 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h74))
				regs_116 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h75))
				regs_117 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h76))
				regs_118 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h77))
				regs_119 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h78))
				regs_120 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h79))
				regs_121 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h7a))
				regs_122 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h7b))
				regs_123 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h7c))
				regs_124 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h7d))
				regs_125 <= io_dst1data_0;
			if (io_wen_0 & (effectiveDst1 == 7'h7e))
				regs_126 <= io_dst1data_0;
			if (io_wen_0 & (&effectiveDst1))
				regs_127 <= io_dst1data_0;
		end
	initial begin : sv2v_autoblock_1
		reg [31:0] _RANDOM [0:127];
	end
	assign io_src1data = io_src1data_0;
	assign io_src2data = io_src2data_0;
endmodule
module TetraNyteCore_Anon (
	io_a,
	io_b,
	io_fn,
	io_out
);
	input [31:0] io_a;
	input [31:0] io_b;
	input [4:0] io_fn;
	output wire [31:0] io_out;
	wire [31:0] io_a_0 = io_a;
	wire [31:0] io_b_0 = io_b;
	wire [4:0] io_fn_0 = io_fn;
	wire [32:0] _GEN = {1'h0, io_a_0};
	wire [32:0] _GEN_0 = {1'h0, io_b_0};
	wire [32:0] _io_out_T = _GEN + _GEN_0;
	wire [31:0] _io_out_T_1 = _io_out_T[31:0];
	wire [32:0] _io_out_T_2 = _GEN - _GEN_0;
	wire [31:0] _io_out_T_3 = _io_out_T_2[31:0];
	wire [31:0] io_out_0 = (io_fn_0 == 5'h00 ? _io_out_T_1 : (io_fn_0 == 5'h01 ? _io_out_T_3 : 32'h00000000));
	assign io_out = io_out_0;
endmodule
module instrMem_1024x32 (
	R0_addr,
	R0_en,
	R0_clk,
	R0_data,
	W0_addr,
	W0_en,
	W0_clk,
	W0_data
);
	input [9:0] R0_addr;
	input R0_en;
	input R0_clk;
	output wire [31:0] R0_data;
	input [9:0] W0_addr;
	input W0_en;
	input W0_clk;
	input [31:0] W0_data;
	reg [31:0] Memory [0:1023];
	reg _R0_en_d0;
	reg [9:0] _R0_addr_d0;
	always @(posedge R0_clk) begin
		_R0_en_d0 <= R0_en;
		_R0_addr_d0 <= R0_addr;
	end
	always @(posedge W0_clk)
		if (W0_en & 1'h1)
			Memory[W0_addr] <= W0_data;
	assign R0_data = (_R0_en_d0 ? Memory[_R0_addr_d0] : 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx);
endmodule
module TetraNyteCore (
	clock,
	reset,
	io_memAddr,
	io_memWdata,
	io_memRdata,
	io_memWe,
	io_instrWriteEnable,
	io_instrWriteAddr,
	io_instrWriteData,
	io_debug
);
	input clock;
	input reset;
	output wire [31:0] io_memAddr;
	output wire [31:0] io_memWdata;
	input [31:0] io_memRdata;
	output wire io_memWe;
	input io_instrWriteEnable;
	input [9:0] io_instrWriteAddr;
	input [31:0] io_instrWriteData;
	input io_debug;
	wire [31:0] io_memRdata_0 = io_memRdata;
	wire io_instrWriteEnable_0 = io_instrWriteEnable;
	wire [9:0] io_instrWriteAddr_0 = io_instrWriteAddr;
	wire [31:0] io_instrWriteData_0 = io_instrWriteData;
	wire io_debug_0 = io_debug;
	wire ifWire_valid = 1'h1;
	wire [1:0] _ifStage_WIRE_threadId = 2'h0;
	wire [1:0] _ifStage_WIRE_1_threadId = 2'h0;
	wire [1:0] _ifStage_WIRE_2_threadId = 2'h0;
	wire [1:0] _ifStage_WIRE_3_threadId = 2'h0;
	wire [1:0] _ifStage_WIRE_4_0_threadId = 2'h0;
	wire [1:0] _ifStage_WIRE_4_1_threadId = 2'h0;
	wire [1:0] _ifStage_WIRE_4_2_threadId = 2'h0;
	wire [1:0] _ifStage_WIRE_4_3_threadId = 2'h0;
	wire [1:0] _decStage_WIRE_threadId = 2'h0;
	wire [1:0] _decStage_WIRE_1_threadId = 2'h0;
	wire [1:0] _decStage_WIRE_2_threadId = 2'h0;
	wire [1:0] _decStage_WIRE_3_threadId = 2'h0;
	wire [1:0] _decStage_WIRE_4_0_threadId = 2'h0;
	wire [1:0] _decStage_WIRE_4_1_threadId = 2'h0;
	wire [1:0] _decStage_WIRE_4_2_threadId = 2'h0;
	wire [1:0] _decStage_WIRE_4_3_threadId = 2'h0;
	wire [1:0] _exStage_WIRE_threadId = 2'h0;
	wire [1:0] _exStage_WIRE_1_threadId = 2'h0;
	wire [1:0] _exStage_WIRE_2_threadId = 2'h0;
	wire [1:0] _exStage_WIRE_3_threadId = 2'h0;
	wire [1:0] _exStage_WIRE_4_0_threadId = 2'h0;
	wire [1:0] _exStage_WIRE_4_1_threadId = 2'h0;
	wire [1:0] _exStage_WIRE_4_2_threadId = 2'h0;
	wire [1:0] _exStage_WIRE_4_3_threadId = 2'h0;
	wire [1:0] _memStage_WIRE_threadId = 2'h0;
	wire [1:0] _memStage_WIRE_1_threadId = 2'h0;
	wire [1:0] _memStage_WIRE_2_threadId = 2'h0;
	wire [1:0] _memStage_WIRE_3_threadId = 2'h0;
	wire [1:0] _memStage_WIRE_4_0_threadId = 2'h0;
	wire [1:0] _memStage_WIRE_4_1_threadId = 2'h0;
	wire [1:0] _memStage_WIRE_4_2_threadId = 2'h0;
	wire [1:0] _memStage_WIRE_4_3_threadId = 2'h0;
	wire [1:0] _ifWire_WIRE_threadId = 2'h0;
	wire [1:0] _decWire_WIRE_threadId = 2'h0;
	wire [1:0] _exWire_WIRE_threadId = 2'h0;
	wire [1:0] _memWire_WIRE_threadId = 2'h0;
	wire _ifStage_WIRE_valid = 1'h0;
	wire _ifStage_WIRE_isALU = 1'h0;
	wire _ifStage_WIRE_isLoad = 1'h0;
	wire _ifStage_WIRE_isStore = 1'h0;
	wire _ifStage_WIRE_isBranch = 1'h0;
	wire _ifStage_WIRE_isJAL = 1'h0;
	wire _ifStage_WIRE_isJALR = 1'h0;
	wire _ifStage_WIRE_isLUI = 1'h0;
	wire _ifStage_WIRE_isAUIPC = 1'h0;
	wire _ifStage_WIRE_isFence = 1'h0;
	wire _ifStage_WIRE_isSystem = 1'h0;
	wire _ifStage_WIRE_1_valid = 1'h0;
	wire _ifStage_WIRE_1_isALU = 1'h0;
	wire _ifStage_WIRE_1_isLoad = 1'h0;
	wire _ifStage_WIRE_1_isStore = 1'h0;
	wire _ifStage_WIRE_1_isBranch = 1'h0;
	wire _ifStage_WIRE_1_isJAL = 1'h0;
	wire _ifStage_WIRE_1_isJALR = 1'h0;
	wire _ifStage_WIRE_1_isLUI = 1'h0;
	wire _ifStage_WIRE_1_isAUIPC = 1'h0;
	wire _ifStage_WIRE_1_isFence = 1'h0;
	wire _ifStage_WIRE_1_isSystem = 1'h0;
	wire _ifStage_WIRE_2_valid = 1'h0;
	wire _ifStage_WIRE_2_isALU = 1'h0;
	wire _ifStage_WIRE_2_isLoad = 1'h0;
	wire _ifStage_WIRE_2_isStore = 1'h0;
	wire _ifStage_WIRE_2_isBranch = 1'h0;
	wire _ifStage_WIRE_2_isJAL = 1'h0;
	wire _ifStage_WIRE_2_isJALR = 1'h0;
	wire _ifStage_WIRE_2_isLUI = 1'h0;
	wire _ifStage_WIRE_2_isAUIPC = 1'h0;
	wire _ifStage_WIRE_2_isFence = 1'h0;
	wire _ifStage_WIRE_2_isSystem = 1'h0;
	wire _ifStage_WIRE_3_valid = 1'h0;
	wire _ifStage_WIRE_3_isALU = 1'h0;
	wire _ifStage_WIRE_3_isLoad = 1'h0;
	wire _ifStage_WIRE_3_isStore = 1'h0;
	wire _ifStage_WIRE_3_isBranch = 1'h0;
	wire _ifStage_WIRE_3_isJAL = 1'h0;
	wire _ifStage_WIRE_3_isJALR = 1'h0;
	wire _ifStage_WIRE_3_isLUI = 1'h0;
	wire _ifStage_WIRE_3_isAUIPC = 1'h0;
	wire _ifStage_WIRE_3_isFence = 1'h0;
	wire _ifStage_WIRE_3_isSystem = 1'h0;
	wire _ifStage_WIRE_4_0_valid = 1'h0;
	wire _ifStage_WIRE_4_0_isALU = 1'h0;
	wire _ifStage_WIRE_4_0_isLoad = 1'h0;
	wire _ifStage_WIRE_4_0_isStore = 1'h0;
	wire _ifStage_WIRE_4_0_isBranch = 1'h0;
	wire _ifStage_WIRE_4_0_isJAL = 1'h0;
	wire _ifStage_WIRE_4_0_isJALR = 1'h0;
	wire _ifStage_WIRE_4_0_isLUI = 1'h0;
	wire _ifStage_WIRE_4_0_isAUIPC = 1'h0;
	wire _ifStage_WIRE_4_0_isFence = 1'h0;
	wire _ifStage_WIRE_4_0_isSystem = 1'h0;
	wire _ifStage_WIRE_4_1_valid = 1'h0;
	wire _ifStage_WIRE_4_1_isALU = 1'h0;
	wire _ifStage_WIRE_4_1_isLoad = 1'h0;
	wire _ifStage_WIRE_4_1_isStore = 1'h0;
	wire _ifStage_WIRE_4_1_isBranch = 1'h0;
	wire _ifStage_WIRE_4_1_isJAL = 1'h0;
	wire _ifStage_WIRE_4_1_isJALR = 1'h0;
	wire _ifStage_WIRE_4_1_isLUI = 1'h0;
	wire _ifStage_WIRE_4_1_isAUIPC = 1'h0;
	wire _ifStage_WIRE_4_1_isFence = 1'h0;
	wire _ifStage_WIRE_4_1_isSystem = 1'h0;
	wire _ifStage_WIRE_4_2_valid = 1'h0;
	wire _ifStage_WIRE_4_2_isALU = 1'h0;
	wire _ifStage_WIRE_4_2_isLoad = 1'h0;
	wire _ifStage_WIRE_4_2_isStore = 1'h0;
	wire _ifStage_WIRE_4_2_isBranch = 1'h0;
	wire _ifStage_WIRE_4_2_isJAL = 1'h0;
	wire _ifStage_WIRE_4_2_isJALR = 1'h0;
	wire _ifStage_WIRE_4_2_isLUI = 1'h0;
	wire _ifStage_WIRE_4_2_isAUIPC = 1'h0;
	wire _ifStage_WIRE_4_2_isFence = 1'h0;
	wire _ifStage_WIRE_4_2_isSystem = 1'h0;
	wire _ifStage_WIRE_4_3_valid = 1'h0;
	wire _ifStage_WIRE_4_3_isALU = 1'h0;
	wire _ifStage_WIRE_4_3_isLoad = 1'h0;
	wire _ifStage_WIRE_4_3_isStore = 1'h0;
	wire _ifStage_WIRE_4_3_isBranch = 1'h0;
	wire _ifStage_WIRE_4_3_isJAL = 1'h0;
	wire _ifStage_WIRE_4_3_isJALR = 1'h0;
	wire _ifStage_WIRE_4_3_isLUI = 1'h0;
	wire _ifStage_WIRE_4_3_isAUIPC = 1'h0;
	wire _ifStage_WIRE_4_3_isFence = 1'h0;
	wire _ifStage_WIRE_4_3_isSystem = 1'h0;
	wire _decStage_WIRE_valid = 1'h0;
	wire _decStage_WIRE_isALU = 1'h0;
	wire _decStage_WIRE_isLoad = 1'h0;
	wire _decStage_WIRE_isStore = 1'h0;
	wire _decStage_WIRE_isBranch = 1'h0;
	wire _decStage_WIRE_isJAL = 1'h0;
	wire _decStage_WIRE_isJALR = 1'h0;
	wire _decStage_WIRE_isLUI = 1'h0;
	wire _decStage_WIRE_isAUIPC = 1'h0;
	wire _decStage_WIRE_isFence = 1'h0;
	wire _decStage_WIRE_isSystem = 1'h0;
	wire _decStage_WIRE_1_valid = 1'h0;
	wire _decStage_WIRE_1_isALU = 1'h0;
	wire _decStage_WIRE_1_isLoad = 1'h0;
	wire _decStage_WIRE_1_isStore = 1'h0;
	wire _decStage_WIRE_1_isBranch = 1'h0;
	wire _decStage_WIRE_1_isJAL = 1'h0;
	wire _decStage_WIRE_1_isJALR = 1'h0;
	wire _decStage_WIRE_1_isLUI = 1'h0;
	wire _decStage_WIRE_1_isAUIPC = 1'h0;
	wire _decStage_WIRE_1_isFence = 1'h0;
	wire _decStage_WIRE_1_isSystem = 1'h0;
	wire _decStage_WIRE_2_valid = 1'h0;
	wire _decStage_WIRE_2_isALU = 1'h0;
	wire _decStage_WIRE_2_isLoad = 1'h0;
	wire _decStage_WIRE_2_isStore = 1'h0;
	wire _decStage_WIRE_2_isBranch = 1'h0;
	wire _decStage_WIRE_2_isJAL = 1'h0;
	wire _decStage_WIRE_2_isJALR = 1'h0;
	wire _decStage_WIRE_2_isLUI = 1'h0;
	wire _decStage_WIRE_2_isAUIPC = 1'h0;
	wire _decStage_WIRE_2_isFence = 1'h0;
	wire _decStage_WIRE_2_isSystem = 1'h0;
	wire _decStage_WIRE_3_valid = 1'h0;
	wire _decStage_WIRE_3_isALU = 1'h0;
	wire _decStage_WIRE_3_isLoad = 1'h0;
	wire _decStage_WIRE_3_isStore = 1'h0;
	wire _decStage_WIRE_3_isBranch = 1'h0;
	wire _decStage_WIRE_3_isJAL = 1'h0;
	wire _decStage_WIRE_3_isJALR = 1'h0;
	wire _decStage_WIRE_3_isLUI = 1'h0;
	wire _decStage_WIRE_3_isAUIPC = 1'h0;
	wire _decStage_WIRE_3_isFence = 1'h0;
	wire _decStage_WIRE_3_isSystem = 1'h0;
	wire _decStage_WIRE_4_0_valid = 1'h0;
	wire _decStage_WIRE_4_0_isALU = 1'h0;
	wire _decStage_WIRE_4_0_isLoad = 1'h0;
	wire _decStage_WIRE_4_0_isStore = 1'h0;
	wire _decStage_WIRE_4_0_isBranch = 1'h0;
	wire _decStage_WIRE_4_0_isJAL = 1'h0;
	wire _decStage_WIRE_4_0_isJALR = 1'h0;
	wire _decStage_WIRE_4_0_isLUI = 1'h0;
	wire _decStage_WIRE_4_0_isAUIPC = 1'h0;
	wire _decStage_WIRE_4_0_isFence = 1'h0;
	wire _decStage_WIRE_4_0_isSystem = 1'h0;
	wire _decStage_WIRE_4_1_valid = 1'h0;
	wire _decStage_WIRE_4_1_isALU = 1'h0;
	wire _decStage_WIRE_4_1_isLoad = 1'h0;
	wire _decStage_WIRE_4_1_isStore = 1'h0;
	wire _decStage_WIRE_4_1_isBranch = 1'h0;
	wire _decStage_WIRE_4_1_isJAL = 1'h0;
	wire _decStage_WIRE_4_1_isJALR = 1'h0;
	wire _decStage_WIRE_4_1_isLUI = 1'h0;
	wire _decStage_WIRE_4_1_isAUIPC = 1'h0;
	wire _decStage_WIRE_4_1_isFence = 1'h0;
	wire _decStage_WIRE_4_1_isSystem = 1'h0;
	wire _decStage_WIRE_4_2_valid = 1'h0;
	wire _decStage_WIRE_4_2_isALU = 1'h0;
	wire _decStage_WIRE_4_2_isLoad = 1'h0;
	wire _decStage_WIRE_4_2_isStore = 1'h0;
	wire _decStage_WIRE_4_2_isBranch = 1'h0;
	wire _decStage_WIRE_4_2_isJAL = 1'h0;
	wire _decStage_WIRE_4_2_isJALR = 1'h0;
	wire _decStage_WIRE_4_2_isLUI = 1'h0;
	wire _decStage_WIRE_4_2_isAUIPC = 1'h0;
	wire _decStage_WIRE_4_2_isFence = 1'h0;
	wire _decStage_WIRE_4_2_isSystem = 1'h0;
	wire _decStage_WIRE_4_3_valid = 1'h0;
	wire _decStage_WIRE_4_3_isALU = 1'h0;
	wire _decStage_WIRE_4_3_isLoad = 1'h0;
	wire _decStage_WIRE_4_3_isStore = 1'h0;
	wire _decStage_WIRE_4_3_isBranch = 1'h0;
	wire _decStage_WIRE_4_3_isJAL = 1'h0;
	wire _decStage_WIRE_4_3_isJALR = 1'h0;
	wire _decStage_WIRE_4_3_isLUI = 1'h0;
	wire _decStage_WIRE_4_3_isAUIPC = 1'h0;
	wire _decStage_WIRE_4_3_isFence = 1'h0;
	wire _decStage_WIRE_4_3_isSystem = 1'h0;
	wire _exStage_WIRE_valid = 1'h0;
	wire _exStage_WIRE_isALU = 1'h0;
	wire _exStage_WIRE_isLoad = 1'h0;
	wire _exStage_WIRE_isStore = 1'h0;
	wire _exStage_WIRE_isBranch = 1'h0;
	wire _exStage_WIRE_isJAL = 1'h0;
	wire _exStage_WIRE_isJALR = 1'h0;
	wire _exStage_WIRE_isLUI = 1'h0;
	wire _exStage_WIRE_isAUIPC = 1'h0;
	wire _exStage_WIRE_isFence = 1'h0;
	wire _exStage_WIRE_isSystem = 1'h0;
	wire _exStage_WIRE_1_valid = 1'h0;
	wire _exStage_WIRE_1_isALU = 1'h0;
	wire _exStage_WIRE_1_isLoad = 1'h0;
	wire _exStage_WIRE_1_isStore = 1'h0;
	wire _exStage_WIRE_1_isBranch = 1'h0;
	wire _exStage_WIRE_1_isJAL = 1'h0;
	wire _exStage_WIRE_1_isJALR = 1'h0;
	wire _exStage_WIRE_1_isLUI = 1'h0;
	wire _exStage_WIRE_1_isAUIPC = 1'h0;
	wire _exStage_WIRE_1_isFence = 1'h0;
	wire _exStage_WIRE_1_isSystem = 1'h0;
	wire _exStage_WIRE_2_valid = 1'h0;
	wire _exStage_WIRE_2_isALU = 1'h0;
	wire _exStage_WIRE_2_isLoad = 1'h0;
	wire _exStage_WIRE_2_isStore = 1'h0;
	wire _exStage_WIRE_2_isBranch = 1'h0;
	wire _exStage_WIRE_2_isJAL = 1'h0;
	wire _exStage_WIRE_2_isJALR = 1'h0;
	wire _exStage_WIRE_2_isLUI = 1'h0;
	wire _exStage_WIRE_2_isAUIPC = 1'h0;
	wire _exStage_WIRE_2_isFence = 1'h0;
	wire _exStage_WIRE_2_isSystem = 1'h0;
	wire _exStage_WIRE_3_valid = 1'h0;
	wire _exStage_WIRE_3_isALU = 1'h0;
	wire _exStage_WIRE_3_isLoad = 1'h0;
	wire _exStage_WIRE_3_isStore = 1'h0;
	wire _exStage_WIRE_3_isBranch = 1'h0;
	wire _exStage_WIRE_3_isJAL = 1'h0;
	wire _exStage_WIRE_3_isJALR = 1'h0;
	wire _exStage_WIRE_3_isLUI = 1'h0;
	wire _exStage_WIRE_3_isAUIPC = 1'h0;
	wire _exStage_WIRE_3_isFence = 1'h0;
	wire _exStage_WIRE_3_isSystem = 1'h0;
	wire _exStage_WIRE_4_0_valid = 1'h0;
	wire _exStage_WIRE_4_0_isALU = 1'h0;
	wire _exStage_WIRE_4_0_isLoad = 1'h0;
	wire _exStage_WIRE_4_0_isStore = 1'h0;
	wire _exStage_WIRE_4_0_isBranch = 1'h0;
	wire _exStage_WIRE_4_0_isJAL = 1'h0;
	wire _exStage_WIRE_4_0_isJALR = 1'h0;
	wire _exStage_WIRE_4_0_isLUI = 1'h0;
	wire _exStage_WIRE_4_0_isAUIPC = 1'h0;
	wire _exStage_WIRE_4_0_isFence = 1'h0;
	wire _exStage_WIRE_4_0_isSystem = 1'h0;
	wire _exStage_WIRE_4_1_valid = 1'h0;
	wire _exStage_WIRE_4_1_isALU = 1'h0;
	wire _exStage_WIRE_4_1_isLoad = 1'h0;
	wire _exStage_WIRE_4_1_isStore = 1'h0;
	wire _exStage_WIRE_4_1_isBranch = 1'h0;
	wire _exStage_WIRE_4_1_isJAL = 1'h0;
	wire _exStage_WIRE_4_1_isJALR = 1'h0;
	wire _exStage_WIRE_4_1_isLUI = 1'h0;
	wire _exStage_WIRE_4_1_isAUIPC = 1'h0;
	wire _exStage_WIRE_4_1_isFence = 1'h0;
	wire _exStage_WIRE_4_1_isSystem = 1'h0;
	wire _exStage_WIRE_4_2_valid = 1'h0;
	wire _exStage_WIRE_4_2_isALU = 1'h0;
	wire _exStage_WIRE_4_2_isLoad = 1'h0;
	wire _exStage_WIRE_4_2_isStore = 1'h0;
	wire _exStage_WIRE_4_2_isBranch = 1'h0;
	wire _exStage_WIRE_4_2_isJAL = 1'h0;
	wire _exStage_WIRE_4_2_isJALR = 1'h0;
	wire _exStage_WIRE_4_2_isLUI = 1'h0;
	wire _exStage_WIRE_4_2_isAUIPC = 1'h0;
	wire _exStage_WIRE_4_2_isFence = 1'h0;
	wire _exStage_WIRE_4_2_isSystem = 1'h0;
	wire _exStage_WIRE_4_3_valid = 1'h0;
	wire _exStage_WIRE_4_3_isALU = 1'h0;
	wire _exStage_WIRE_4_3_isLoad = 1'h0;
	wire _exStage_WIRE_4_3_isStore = 1'h0;
	wire _exStage_WIRE_4_3_isBranch = 1'h0;
	wire _exStage_WIRE_4_3_isJAL = 1'h0;
	wire _exStage_WIRE_4_3_isJALR = 1'h0;
	wire _exStage_WIRE_4_3_isLUI = 1'h0;
	wire _exStage_WIRE_4_3_isAUIPC = 1'h0;
	wire _exStage_WIRE_4_3_isFence = 1'h0;
	wire _exStage_WIRE_4_3_isSystem = 1'h0;
	wire _memStage_WIRE_valid = 1'h0;
	wire _memStage_WIRE_isALU = 1'h0;
	wire _memStage_WIRE_isLoad = 1'h0;
	wire _memStage_WIRE_isStore = 1'h0;
	wire _memStage_WIRE_isBranch = 1'h0;
	wire _memStage_WIRE_isJAL = 1'h0;
	wire _memStage_WIRE_isJALR = 1'h0;
	wire _memStage_WIRE_isLUI = 1'h0;
	wire _memStage_WIRE_isAUIPC = 1'h0;
	wire _memStage_WIRE_isFence = 1'h0;
	wire _memStage_WIRE_isSystem = 1'h0;
	wire _memStage_WIRE_1_valid = 1'h0;
	wire _memStage_WIRE_1_isALU = 1'h0;
	wire _memStage_WIRE_1_isLoad = 1'h0;
	wire _memStage_WIRE_1_isStore = 1'h0;
	wire _memStage_WIRE_1_isBranch = 1'h0;
	wire _memStage_WIRE_1_isJAL = 1'h0;
	wire _memStage_WIRE_1_isJALR = 1'h0;
	wire _memStage_WIRE_1_isLUI = 1'h0;
	wire _memStage_WIRE_1_isAUIPC = 1'h0;
	wire _memStage_WIRE_1_isFence = 1'h0;
	wire _memStage_WIRE_1_isSystem = 1'h0;
	wire _memStage_WIRE_2_valid = 1'h0;
	wire _memStage_WIRE_2_isALU = 1'h0;
	wire _memStage_WIRE_2_isLoad = 1'h0;
	wire _memStage_WIRE_2_isStore = 1'h0;
	wire _memStage_WIRE_2_isBranch = 1'h0;
	wire _memStage_WIRE_2_isJAL = 1'h0;
	wire _memStage_WIRE_2_isJALR = 1'h0;
	wire _memStage_WIRE_2_isLUI = 1'h0;
	wire _memStage_WIRE_2_isAUIPC = 1'h0;
	wire _memStage_WIRE_2_isFence = 1'h0;
	wire _memStage_WIRE_2_isSystem = 1'h0;
	wire _memStage_WIRE_3_valid = 1'h0;
	wire _memStage_WIRE_3_isALU = 1'h0;
	wire _memStage_WIRE_3_isLoad = 1'h0;
	wire _memStage_WIRE_3_isStore = 1'h0;
	wire _memStage_WIRE_3_isBranch = 1'h0;
	wire _memStage_WIRE_3_isJAL = 1'h0;
	wire _memStage_WIRE_3_isJALR = 1'h0;
	wire _memStage_WIRE_3_isLUI = 1'h0;
	wire _memStage_WIRE_3_isAUIPC = 1'h0;
	wire _memStage_WIRE_3_isFence = 1'h0;
	wire _memStage_WIRE_3_isSystem = 1'h0;
	wire _memStage_WIRE_4_0_valid = 1'h0;
	wire _memStage_WIRE_4_0_isALU = 1'h0;
	wire _memStage_WIRE_4_0_isLoad = 1'h0;
	wire _memStage_WIRE_4_0_isStore = 1'h0;
	wire _memStage_WIRE_4_0_isBranch = 1'h0;
	wire _memStage_WIRE_4_0_isJAL = 1'h0;
	wire _memStage_WIRE_4_0_isJALR = 1'h0;
	wire _memStage_WIRE_4_0_isLUI = 1'h0;
	wire _memStage_WIRE_4_0_isAUIPC = 1'h0;
	wire _memStage_WIRE_4_0_isFence = 1'h0;
	wire _memStage_WIRE_4_0_isSystem = 1'h0;
	wire _memStage_WIRE_4_1_valid = 1'h0;
	wire _memStage_WIRE_4_1_isALU = 1'h0;
	wire _memStage_WIRE_4_1_isLoad = 1'h0;
	wire _memStage_WIRE_4_1_isStore = 1'h0;
	wire _memStage_WIRE_4_1_isBranch = 1'h0;
	wire _memStage_WIRE_4_1_isJAL = 1'h0;
	wire _memStage_WIRE_4_1_isJALR = 1'h0;
	wire _memStage_WIRE_4_1_isLUI = 1'h0;
	wire _memStage_WIRE_4_1_isAUIPC = 1'h0;
	wire _memStage_WIRE_4_1_isFence = 1'h0;
	wire _memStage_WIRE_4_1_isSystem = 1'h0;
	wire _memStage_WIRE_4_2_valid = 1'h0;
	wire _memStage_WIRE_4_2_isALU = 1'h0;
	wire _memStage_WIRE_4_2_isLoad = 1'h0;
	wire _memStage_WIRE_4_2_isStore = 1'h0;
	wire _memStage_WIRE_4_2_isBranch = 1'h0;
	wire _memStage_WIRE_4_2_isJAL = 1'h0;
	wire _memStage_WIRE_4_2_isJALR = 1'h0;
	wire _memStage_WIRE_4_2_isLUI = 1'h0;
	wire _memStage_WIRE_4_2_isAUIPC = 1'h0;
	wire _memStage_WIRE_4_2_isFence = 1'h0;
	wire _memStage_WIRE_4_2_isSystem = 1'h0;
	wire _memStage_WIRE_4_3_valid = 1'h0;
	wire _memStage_WIRE_4_3_isALU = 1'h0;
	wire _memStage_WIRE_4_3_isLoad = 1'h0;
	wire _memStage_WIRE_4_3_isStore = 1'h0;
	wire _memStage_WIRE_4_3_isBranch = 1'h0;
	wire _memStage_WIRE_4_3_isJAL = 1'h0;
	wire _memStage_WIRE_4_3_isJALR = 1'h0;
	wire _memStage_WIRE_4_3_isLUI = 1'h0;
	wire _memStage_WIRE_4_3_isAUIPC = 1'h0;
	wire _memStage_WIRE_4_3_isFence = 1'h0;
	wire _memStage_WIRE_4_3_isSystem = 1'h0;
	wire _ifWire_WIRE_valid = 1'h0;
	wire _ifWire_WIRE_isALU = 1'h0;
	wire _ifWire_WIRE_isLoad = 1'h0;
	wire _ifWire_WIRE_isStore = 1'h0;
	wire _ifWire_WIRE_isBranch = 1'h0;
	wire _ifWire_WIRE_isJAL = 1'h0;
	wire _ifWire_WIRE_isJALR = 1'h0;
	wire _ifWire_WIRE_isLUI = 1'h0;
	wire _ifWire_WIRE_isAUIPC = 1'h0;
	wire _ifWire_WIRE_isFence = 1'h0;
	wire _ifWire_WIRE_isSystem = 1'h0;
	wire ifWire_isALU = 1'h0;
	wire ifWire_isLoad = 1'h0;
	wire ifWire_isStore = 1'h0;
	wire ifWire_isBranch = 1'h0;
	wire ifWire_isJAL = 1'h0;
	wire ifWire_isJALR = 1'h0;
	wire ifWire_isLUI = 1'h0;
	wire ifWire_isAUIPC = 1'h0;
	wire ifWire_isFence = 1'h0;
	wire ifWire_isSystem = 1'h0;
	wire _decWire_WIRE_valid = 1'h0;
	wire _decWire_WIRE_isALU = 1'h0;
	wire _decWire_WIRE_isLoad = 1'h0;
	wire _decWire_WIRE_isStore = 1'h0;
	wire _decWire_WIRE_isBranch = 1'h0;
	wire _decWire_WIRE_isJAL = 1'h0;
	wire _decWire_WIRE_isJALR = 1'h0;
	wire _decWire_WIRE_isLUI = 1'h0;
	wire _decWire_WIRE_isAUIPC = 1'h0;
	wire _decWire_WIRE_isFence = 1'h0;
	wire _decWire_WIRE_isSystem = 1'h0;
	wire _exWire_WIRE_valid = 1'h0;
	wire _exWire_WIRE_isALU = 1'h0;
	wire _exWire_WIRE_isLoad = 1'h0;
	wire _exWire_WIRE_isStore = 1'h0;
	wire _exWire_WIRE_isBranch = 1'h0;
	wire _exWire_WIRE_isJAL = 1'h0;
	wire _exWire_WIRE_isJALR = 1'h0;
	wire _exWire_WIRE_isLUI = 1'h0;
	wire _exWire_WIRE_isAUIPC = 1'h0;
	wire _exWire_WIRE_isFence = 1'h0;
	wire _exWire_WIRE_isSystem = 1'h0;
	wire _memWire_WIRE_valid = 1'h0;
	wire _memWire_WIRE_isALU = 1'h0;
	wire _memWire_WIRE_isLoad = 1'h0;
	wire _memWire_WIRE_isStore = 1'h0;
	wire _memWire_WIRE_isBranch = 1'h0;
	wire _memWire_WIRE_isJAL = 1'h0;
	wire _memWire_WIRE_isJALR = 1'h0;
	wire _memWire_WIRE_isLUI = 1'h0;
	wire _memWire_WIRE_isAUIPC = 1'h0;
	wire _memWire_WIRE_isFence = 1'h0;
	wire _memWire_WIRE_isSystem = 1'h0;
	wire [4:0] _ifStage_WIRE_aluOp = 5'h00;
	wire [4:0] _ifStage_WIRE_rs1 = 5'h00;
	wire [4:0] _ifStage_WIRE_rs2 = 5'h00;
	wire [4:0] _ifStage_WIRE_rd = 5'h00;
	wire [4:0] _ifStage_WIRE_1_aluOp = 5'h00;
	wire [4:0] _ifStage_WIRE_1_rs1 = 5'h00;
	wire [4:0] _ifStage_WIRE_1_rs2 = 5'h00;
	wire [4:0] _ifStage_WIRE_1_rd = 5'h00;
	wire [4:0] _ifStage_WIRE_2_aluOp = 5'h00;
	wire [4:0] _ifStage_WIRE_2_rs1 = 5'h00;
	wire [4:0] _ifStage_WIRE_2_rs2 = 5'h00;
	wire [4:0] _ifStage_WIRE_2_rd = 5'h00;
	wire [4:0] _ifStage_WIRE_3_aluOp = 5'h00;
	wire [4:0] _ifStage_WIRE_3_rs1 = 5'h00;
	wire [4:0] _ifStage_WIRE_3_rs2 = 5'h00;
	wire [4:0] _ifStage_WIRE_3_rd = 5'h00;
	wire [4:0] _ifStage_WIRE_4_0_aluOp = 5'h00;
	wire [4:0] _ifStage_WIRE_4_0_rs1 = 5'h00;
	wire [4:0] _ifStage_WIRE_4_0_rs2 = 5'h00;
	wire [4:0] _ifStage_WIRE_4_0_rd = 5'h00;
	wire [4:0] _ifStage_WIRE_4_1_aluOp = 5'h00;
	wire [4:0] _ifStage_WIRE_4_1_rs1 = 5'h00;
	wire [4:0] _ifStage_WIRE_4_1_rs2 = 5'h00;
	wire [4:0] _ifStage_WIRE_4_1_rd = 5'h00;
	wire [4:0] _ifStage_WIRE_4_2_aluOp = 5'h00;
	wire [4:0] _ifStage_WIRE_4_2_rs1 = 5'h00;
	wire [4:0] _ifStage_WIRE_4_2_rs2 = 5'h00;
	wire [4:0] _ifStage_WIRE_4_2_rd = 5'h00;
	wire [4:0] _ifStage_WIRE_4_3_aluOp = 5'h00;
	wire [4:0] _ifStage_WIRE_4_3_rs1 = 5'h00;
	wire [4:0] _ifStage_WIRE_4_3_rs2 = 5'h00;
	wire [4:0] _ifStage_WIRE_4_3_rd = 5'h00;
	wire [4:0] _decStage_WIRE_aluOp = 5'h00;
	wire [4:0] _decStage_WIRE_rs1 = 5'h00;
	wire [4:0] _decStage_WIRE_rs2 = 5'h00;
	wire [4:0] _decStage_WIRE_rd = 5'h00;
	wire [4:0] _decStage_WIRE_1_aluOp = 5'h00;
	wire [4:0] _decStage_WIRE_1_rs1 = 5'h00;
	wire [4:0] _decStage_WIRE_1_rs2 = 5'h00;
	wire [4:0] _decStage_WIRE_1_rd = 5'h00;
	wire [4:0] _decStage_WIRE_2_aluOp = 5'h00;
	wire [4:0] _decStage_WIRE_2_rs1 = 5'h00;
	wire [4:0] _decStage_WIRE_2_rs2 = 5'h00;
	wire [4:0] _decStage_WIRE_2_rd = 5'h00;
	wire [4:0] _decStage_WIRE_3_aluOp = 5'h00;
	wire [4:0] _decStage_WIRE_3_rs1 = 5'h00;
	wire [4:0] _decStage_WIRE_3_rs2 = 5'h00;
	wire [4:0] _decStage_WIRE_3_rd = 5'h00;
	wire [4:0] _decStage_WIRE_4_0_aluOp = 5'h00;
	wire [4:0] _decStage_WIRE_4_0_rs1 = 5'h00;
	wire [4:0] _decStage_WIRE_4_0_rs2 = 5'h00;
	wire [4:0] _decStage_WIRE_4_0_rd = 5'h00;
	wire [4:0] _decStage_WIRE_4_1_aluOp = 5'h00;
	wire [4:0] _decStage_WIRE_4_1_rs1 = 5'h00;
	wire [4:0] _decStage_WIRE_4_1_rs2 = 5'h00;
	wire [4:0] _decStage_WIRE_4_1_rd = 5'h00;
	wire [4:0] _decStage_WIRE_4_2_aluOp = 5'h00;
	wire [4:0] _decStage_WIRE_4_2_rs1 = 5'h00;
	wire [4:0] _decStage_WIRE_4_2_rs2 = 5'h00;
	wire [4:0] _decStage_WIRE_4_2_rd = 5'h00;
	wire [4:0] _decStage_WIRE_4_3_aluOp = 5'h00;
	wire [4:0] _decStage_WIRE_4_3_rs1 = 5'h00;
	wire [4:0] _decStage_WIRE_4_3_rs2 = 5'h00;
	wire [4:0] _decStage_WIRE_4_3_rd = 5'h00;
	wire [4:0] _exStage_WIRE_aluOp = 5'h00;
	wire [4:0] _exStage_WIRE_rs1 = 5'h00;
	wire [4:0] _exStage_WIRE_rs2 = 5'h00;
	wire [4:0] _exStage_WIRE_rd = 5'h00;
	wire [4:0] _exStage_WIRE_1_aluOp = 5'h00;
	wire [4:0] _exStage_WIRE_1_rs1 = 5'h00;
	wire [4:0] _exStage_WIRE_1_rs2 = 5'h00;
	wire [4:0] _exStage_WIRE_1_rd = 5'h00;
	wire [4:0] _exStage_WIRE_2_aluOp = 5'h00;
	wire [4:0] _exStage_WIRE_2_rs1 = 5'h00;
	wire [4:0] _exStage_WIRE_2_rs2 = 5'h00;
	wire [4:0] _exStage_WIRE_2_rd = 5'h00;
	wire [4:0] _exStage_WIRE_3_aluOp = 5'h00;
	wire [4:0] _exStage_WIRE_3_rs1 = 5'h00;
	wire [4:0] _exStage_WIRE_3_rs2 = 5'h00;
	wire [4:0] _exStage_WIRE_3_rd = 5'h00;
	wire [4:0] _exStage_WIRE_4_0_aluOp = 5'h00;
	wire [4:0] _exStage_WIRE_4_0_rs1 = 5'h00;
	wire [4:0] _exStage_WIRE_4_0_rs2 = 5'h00;
	wire [4:0] _exStage_WIRE_4_0_rd = 5'h00;
	wire [4:0] _exStage_WIRE_4_1_aluOp = 5'h00;
	wire [4:0] _exStage_WIRE_4_1_rs1 = 5'h00;
	wire [4:0] _exStage_WIRE_4_1_rs2 = 5'h00;
	wire [4:0] _exStage_WIRE_4_1_rd = 5'h00;
	wire [4:0] _exStage_WIRE_4_2_aluOp = 5'h00;
	wire [4:0] _exStage_WIRE_4_2_rs1 = 5'h00;
	wire [4:0] _exStage_WIRE_4_2_rs2 = 5'h00;
	wire [4:0] _exStage_WIRE_4_2_rd = 5'h00;
	wire [4:0] _exStage_WIRE_4_3_aluOp = 5'h00;
	wire [4:0] _exStage_WIRE_4_3_rs1 = 5'h00;
	wire [4:0] _exStage_WIRE_4_3_rs2 = 5'h00;
	wire [4:0] _exStage_WIRE_4_3_rd = 5'h00;
	wire [4:0] _memStage_WIRE_aluOp = 5'h00;
	wire [4:0] _memStage_WIRE_rs1 = 5'h00;
	wire [4:0] _memStage_WIRE_rs2 = 5'h00;
	wire [4:0] _memStage_WIRE_rd = 5'h00;
	wire [4:0] _memStage_WIRE_1_aluOp = 5'h00;
	wire [4:0] _memStage_WIRE_1_rs1 = 5'h00;
	wire [4:0] _memStage_WIRE_1_rs2 = 5'h00;
	wire [4:0] _memStage_WIRE_1_rd = 5'h00;
	wire [4:0] _memStage_WIRE_2_aluOp = 5'h00;
	wire [4:0] _memStage_WIRE_2_rs1 = 5'h00;
	wire [4:0] _memStage_WIRE_2_rs2 = 5'h00;
	wire [4:0] _memStage_WIRE_2_rd = 5'h00;
	wire [4:0] _memStage_WIRE_3_aluOp = 5'h00;
	wire [4:0] _memStage_WIRE_3_rs1 = 5'h00;
	wire [4:0] _memStage_WIRE_3_rs2 = 5'h00;
	wire [4:0] _memStage_WIRE_3_rd = 5'h00;
	wire [4:0] _memStage_WIRE_4_0_aluOp = 5'h00;
	wire [4:0] _memStage_WIRE_4_0_rs1 = 5'h00;
	wire [4:0] _memStage_WIRE_4_0_rs2 = 5'h00;
	wire [4:0] _memStage_WIRE_4_0_rd = 5'h00;
	wire [4:0] _memStage_WIRE_4_1_aluOp = 5'h00;
	wire [4:0] _memStage_WIRE_4_1_rs1 = 5'h00;
	wire [4:0] _memStage_WIRE_4_1_rs2 = 5'h00;
	wire [4:0] _memStage_WIRE_4_1_rd = 5'h00;
	wire [4:0] _memStage_WIRE_4_2_aluOp = 5'h00;
	wire [4:0] _memStage_WIRE_4_2_rs1 = 5'h00;
	wire [4:0] _memStage_WIRE_4_2_rs2 = 5'h00;
	wire [4:0] _memStage_WIRE_4_2_rd = 5'h00;
	wire [4:0] _memStage_WIRE_4_3_aluOp = 5'h00;
	wire [4:0] _memStage_WIRE_4_3_rs1 = 5'h00;
	wire [4:0] _memStage_WIRE_4_3_rs2 = 5'h00;
	wire [4:0] _memStage_WIRE_4_3_rd = 5'h00;
	wire [4:0] _ifWire_WIRE_aluOp = 5'h00;
	wire [4:0] _ifWire_WIRE_rs1 = 5'h00;
	wire [4:0] _ifWire_WIRE_rs2 = 5'h00;
	wire [4:0] _ifWire_WIRE_rd = 5'h00;
	wire [4:0] ifWire_aluOp = 5'h00;
	wire [4:0] ifWire_rs1 = 5'h00;
	wire [4:0] ifWire_rs2 = 5'h00;
	wire [4:0] ifWire_rd = 5'h00;
	wire [4:0] _decWire_WIRE_aluOp = 5'h00;
	wire [4:0] _decWire_WIRE_rs1 = 5'h00;
	wire [4:0] _decWire_WIRE_rs2 = 5'h00;
	wire [4:0] _decWire_WIRE_rd = 5'h00;
	wire [4:0] _exWire_WIRE_aluOp = 5'h00;
	wire [4:0] _exWire_WIRE_rs1 = 5'h00;
	wire [4:0] _exWire_WIRE_rs2 = 5'h00;
	wire [4:0] _exWire_WIRE_rd = 5'h00;
	wire [4:0] _memWire_WIRE_aluOp = 5'h00;
	wire [4:0] _memWire_WIRE_rs1 = 5'h00;
	wire [4:0] _memWire_WIRE_rs2 = 5'h00;
	wire [4:0] _memWire_WIRE_rd = 5'h00;
	wire [31:0] _pcRegs_WIRE_0 = 32'h00000000;
	wire [31:0] _pcRegs_WIRE_1 = 32'h00000000;
	wire [31:0] _pcRegs_WIRE_2 = 32'h00000000;
	wire [31:0] _pcRegs_WIRE_3 = 32'h00000000;
	wire [31:0] _ifStage_WIRE_pc = 32'h00000000;
	wire [31:0] _ifStage_WIRE_instr = 32'h00000000;
	wire [31:0] _ifStage_WIRE_imm = 32'h00000000;
	wire [31:0] _ifStage_WIRE_rs1Data = 32'h00000000;
	wire [31:0] _ifStage_WIRE_rs2Data = 32'h00000000;
	wire [31:0] _ifStage_WIRE_memAddr = 32'h00000000;
	wire [31:0] _ifStage_WIRE_memWdata = 32'h00000000;
	wire [31:0] _ifStage_WIRE_memRdata = 32'h00000000;
	wire [31:0] _ifStage_WIRE_aluResult = 32'h00000000;
	wire [31:0] _ifStage_WIRE_1_pc = 32'h00000000;
	wire [31:0] _ifStage_WIRE_1_instr = 32'h00000000;
	wire [31:0] _ifStage_WIRE_1_imm = 32'h00000000;
	wire [31:0] _ifStage_WIRE_1_rs1Data = 32'h00000000;
	wire [31:0] _ifStage_WIRE_1_rs2Data = 32'h00000000;
	wire [31:0] _ifStage_WIRE_1_memAddr = 32'h00000000;
	wire [31:0] _ifStage_WIRE_1_memWdata = 32'h00000000;
	wire [31:0] _ifStage_WIRE_1_memRdata = 32'h00000000;
	wire [31:0] _ifStage_WIRE_1_aluResult = 32'h00000000;
	wire [31:0] _ifStage_WIRE_2_pc = 32'h00000000;
	wire [31:0] _ifStage_WIRE_2_instr = 32'h00000000;
	wire [31:0] _ifStage_WIRE_2_imm = 32'h00000000;
	wire [31:0] _ifStage_WIRE_2_rs1Data = 32'h00000000;
	wire [31:0] _ifStage_WIRE_2_rs2Data = 32'h00000000;
	wire [31:0] _ifStage_WIRE_2_memAddr = 32'h00000000;
	wire [31:0] _ifStage_WIRE_2_memWdata = 32'h00000000;
	wire [31:0] _ifStage_WIRE_2_memRdata = 32'h00000000;
	wire [31:0] _ifStage_WIRE_2_aluResult = 32'h00000000;
	wire [31:0] _ifStage_WIRE_3_pc = 32'h00000000;
	wire [31:0] _ifStage_WIRE_3_instr = 32'h00000000;
	wire [31:0] _ifStage_WIRE_3_imm = 32'h00000000;
	wire [31:0] _ifStage_WIRE_3_rs1Data = 32'h00000000;
	wire [31:0] _ifStage_WIRE_3_rs2Data = 32'h00000000;
	wire [31:0] _ifStage_WIRE_3_memAddr = 32'h00000000;
	wire [31:0] _ifStage_WIRE_3_memWdata = 32'h00000000;
	wire [31:0] _ifStage_WIRE_3_memRdata = 32'h00000000;
	wire [31:0] _ifStage_WIRE_3_aluResult = 32'h00000000;
	wire [31:0] _ifStage_WIRE_4_0_pc = 32'h00000000;
	wire [31:0] _ifStage_WIRE_4_0_instr = 32'h00000000;
	wire [31:0] _ifStage_WIRE_4_0_imm = 32'h00000000;
	wire [31:0] _ifStage_WIRE_4_0_rs1Data = 32'h00000000;
	wire [31:0] _ifStage_WIRE_4_0_rs2Data = 32'h00000000;
	wire [31:0] _ifStage_WIRE_4_0_memAddr = 32'h00000000;
	wire [31:0] _ifStage_WIRE_4_0_memWdata = 32'h00000000;
	wire [31:0] _ifStage_WIRE_4_0_memRdata = 32'h00000000;
	wire [31:0] _ifStage_WIRE_4_0_aluResult = 32'h00000000;
	wire [31:0] _ifStage_WIRE_4_1_pc = 32'h00000000;
	wire [31:0] _ifStage_WIRE_4_1_instr = 32'h00000000;
	wire [31:0] _ifStage_WIRE_4_1_imm = 32'h00000000;
	wire [31:0] _ifStage_WIRE_4_1_rs1Data = 32'h00000000;
	wire [31:0] _ifStage_WIRE_4_1_rs2Data = 32'h00000000;
	wire [31:0] _ifStage_WIRE_4_1_memAddr = 32'h00000000;
	wire [31:0] _ifStage_WIRE_4_1_memWdata = 32'h00000000;
	wire [31:0] _ifStage_WIRE_4_1_memRdata = 32'h00000000;
	wire [31:0] _ifStage_WIRE_4_1_aluResult = 32'h00000000;
	wire [31:0] _ifStage_WIRE_4_2_pc = 32'h00000000;
	wire [31:0] _ifStage_WIRE_4_2_instr = 32'h00000000;
	wire [31:0] _ifStage_WIRE_4_2_imm = 32'h00000000;
	wire [31:0] _ifStage_WIRE_4_2_rs1Data = 32'h00000000;
	wire [31:0] _ifStage_WIRE_4_2_rs2Data = 32'h00000000;
	wire [31:0] _ifStage_WIRE_4_2_memAddr = 32'h00000000;
	wire [31:0] _ifStage_WIRE_4_2_memWdata = 32'h00000000;
	wire [31:0] _ifStage_WIRE_4_2_memRdata = 32'h00000000;
	wire [31:0] _ifStage_WIRE_4_2_aluResult = 32'h00000000;
	wire [31:0] _ifStage_WIRE_4_3_pc = 32'h00000000;
	wire [31:0] _ifStage_WIRE_4_3_instr = 32'h00000000;
	wire [31:0] _ifStage_WIRE_4_3_imm = 32'h00000000;
	wire [31:0] _ifStage_WIRE_4_3_rs1Data = 32'h00000000;
	wire [31:0] _ifStage_WIRE_4_3_rs2Data = 32'h00000000;
	wire [31:0] _ifStage_WIRE_4_3_memAddr = 32'h00000000;
	wire [31:0] _ifStage_WIRE_4_3_memWdata = 32'h00000000;
	wire [31:0] _ifStage_WIRE_4_3_memRdata = 32'h00000000;
	wire [31:0] _ifStage_WIRE_4_3_aluResult = 32'h00000000;
	wire [31:0] _decStage_WIRE_pc = 32'h00000000;
	wire [31:0] _decStage_WIRE_instr = 32'h00000000;
	wire [31:0] _decStage_WIRE_imm = 32'h00000000;
	wire [31:0] _decStage_WIRE_rs1Data = 32'h00000000;
	wire [31:0] _decStage_WIRE_rs2Data = 32'h00000000;
	wire [31:0] _decStage_WIRE_memAddr = 32'h00000000;
	wire [31:0] _decStage_WIRE_memWdata = 32'h00000000;
	wire [31:0] _decStage_WIRE_memRdata = 32'h00000000;
	wire [31:0] _decStage_WIRE_aluResult = 32'h00000000;
	wire [31:0] _decStage_WIRE_1_pc = 32'h00000000;
	wire [31:0] _decStage_WIRE_1_instr = 32'h00000000;
	wire [31:0] _decStage_WIRE_1_imm = 32'h00000000;
	wire [31:0] _decStage_WIRE_1_rs1Data = 32'h00000000;
	wire [31:0] _decStage_WIRE_1_rs2Data = 32'h00000000;
	wire [31:0] _decStage_WIRE_1_memAddr = 32'h00000000;
	wire [31:0] _decStage_WIRE_1_memWdata = 32'h00000000;
	wire [31:0] _decStage_WIRE_1_memRdata = 32'h00000000;
	wire [31:0] _decStage_WIRE_1_aluResult = 32'h00000000;
	wire [31:0] _decStage_WIRE_2_pc = 32'h00000000;
	wire [31:0] _decStage_WIRE_2_instr = 32'h00000000;
	wire [31:0] _decStage_WIRE_2_imm = 32'h00000000;
	wire [31:0] _decStage_WIRE_2_rs1Data = 32'h00000000;
	wire [31:0] _decStage_WIRE_2_rs2Data = 32'h00000000;
	wire [31:0] _decStage_WIRE_2_memAddr = 32'h00000000;
	wire [31:0] _decStage_WIRE_2_memWdata = 32'h00000000;
	wire [31:0] _decStage_WIRE_2_memRdata = 32'h00000000;
	wire [31:0] _decStage_WIRE_2_aluResult = 32'h00000000;
	wire [31:0] _decStage_WIRE_3_pc = 32'h00000000;
	wire [31:0] _decStage_WIRE_3_instr = 32'h00000000;
	wire [31:0] _decStage_WIRE_3_imm = 32'h00000000;
	wire [31:0] _decStage_WIRE_3_rs1Data = 32'h00000000;
	wire [31:0] _decStage_WIRE_3_rs2Data = 32'h00000000;
	wire [31:0] _decStage_WIRE_3_memAddr = 32'h00000000;
	wire [31:0] _decStage_WIRE_3_memWdata = 32'h00000000;
	wire [31:0] _decStage_WIRE_3_memRdata = 32'h00000000;
	wire [31:0] _decStage_WIRE_3_aluResult = 32'h00000000;
	wire [31:0] _decStage_WIRE_4_0_pc = 32'h00000000;
	wire [31:0] _decStage_WIRE_4_0_instr = 32'h00000000;
	wire [31:0] _decStage_WIRE_4_0_imm = 32'h00000000;
	wire [31:0] _decStage_WIRE_4_0_rs1Data = 32'h00000000;
	wire [31:0] _decStage_WIRE_4_0_rs2Data = 32'h00000000;
	wire [31:0] _decStage_WIRE_4_0_memAddr = 32'h00000000;
	wire [31:0] _decStage_WIRE_4_0_memWdata = 32'h00000000;
	wire [31:0] _decStage_WIRE_4_0_memRdata = 32'h00000000;
	wire [31:0] _decStage_WIRE_4_0_aluResult = 32'h00000000;
	wire [31:0] _decStage_WIRE_4_1_pc = 32'h00000000;
	wire [31:0] _decStage_WIRE_4_1_instr = 32'h00000000;
	wire [31:0] _decStage_WIRE_4_1_imm = 32'h00000000;
	wire [31:0] _decStage_WIRE_4_1_rs1Data = 32'h00000000;
	wire [31:0] _decStage_WIRE_4_1_rs2Data = 32'h00000000;
	wire [31:0] _decStage_WIRE_4_1_memAddr = 32'h00000000;
	wire [31:0] _decStage_WIRE_4_1_memWdata = 32'h00000000;
	wire [31:0] _decStage_WIRE_4_1_memRdata = 32'h00000000;
	wire [31:0] _decStage_WIRE_4_1_aluResult = 32'h00000000;
	wire [31:0] _decStage_WIRE_4_2_pc = 32'h00000000;
	wire [31:0] _decStage_WIRE_4_2_instr = 32'h00000000;
	wire [31:0] _decStage_WIRE_4_2_imm = 32'h00000000;
	wire [31:0] _decStage_WIRE_4_2_rs1Data = 32'h00000000;
	wire [31:0] _decStage_WIRE_4_2_rs2Data = 32'h00000000;
	wire [31:0] _decStage_WIRE_4_2_memAddr = 32'h00000000;
	wire [31:0] _decStage_WIRE_4_2_memWdata = 32'h00000000;
	wire [31:0] _decStage_WIRE_4_2_memRdata = 32'h00000000;
	wire [31:0] _decStage_WIRE_4_2_aluResult = 32'h00000000;
	wire [31:0] _decStage_WIRE_4_3_pc = 32'h00000000;
	wire [31:0] _decStage_WIRE_4_3_instr = 32'h00000000;
	wire [31:0] _decStage_WIRE_4_3_imm = 32'h00000000;
	wire [31:0] _decStage_WIRE_4_3_rs1Data = 32'h00000000;
	wire [31:0] _decStage_WIRE_4_3_rs2Data = 32'h00000000;
	wire [31:0] _decStage_WIRE_4_3_memAddr = 32'h00000000;
	wire [31:0] _decStage_WIRE_4_3_memWdata = 32'h00000000;
	wire [31:0] _decStage_WIRE_4_3_memRdata = 32'h00000000;
	wire [31:0] _decStage_WIRE_4_3_aluResult = 32'h00000000;
	wire [31:0] _exStage_WIRE_pc = 32'h00000000;
	wire [31:0] _exStage_WIRE_instr = 32'h00000000;
	wire [31:0] _exStage_WIRE_imm = 32'h00000000;
	wire [31:0] _exStage_WIRE_rs1Data = 32'h00000000;
	wire [31:0] _exStage_WIRE_rs2Data = 32'h00000000;
	wire [31:0] _exStage_WIRE_memAddr = 32'h00000000;
	wire [31:0] _exStage_WIRE_memWdata = 32'h00000000;
	wire [31:0] _exStage_WIRE_memRdata = 32'h00000000;
	wire [31:0] _exStage_WIRE_aluResult = 32'h00000000;
	wire [31:0] _exStage_WIRE_1_pc = 32'h00000000;
	wire [31:0] _exStage_WIRE_1_instr = 32'h00000000;
	wire [31:0] _exStage_WIRE_1_imm = 32'h00000000;
	wire [31:0] _exStage_WIRE_1_rs1Data = 32'h00000000;
	wire [31:0] _exStage_WIRE_1_rs2Data = 32'h00000000;
	wire [31:0] _exStage_WIRE_1_memAddr = 32'h00000000;
	wire [31:0] _exStage_WIRE_1_memWdata = 32'h00000000;
	wire [31:0] _exStage_WIRE_1_memRdata = 32'h00000000;
	wire [31:0] _exStage_WIRE_1_aluResult = 32'h00000000;
	wire [31:0] _exStage_WIRE_2_pc = 32'h00000000;
	wire [31:0] _exStage_WIRE_2_instr = 32'h00000000;
	wire [31:0] _exStage_WIRE_2_imm = 32'h00000000;
	wire [31:0] _exStage_WIRE_2_rs1Data = 32'h00000000;
	wire [31:0] _exStage_WIRE_2_rs2Data = 32'h00000000;
	wire [31:0] _exStage_WIRE_2_memAddr = 32'h00000000;
	wire [31:0] _exStage_WIRE_2_memWdata = 32'h00000000;
	wire [31:0] _exStage_WIRE_2_memRdata = 32'h00000000;
	wire [31:0] _exStage_WIRE_2_aluResult = 32'h00000000;
	wire [31:0] _exStage_WIRE_3_pc = 32'h00000000;
	wire [31:0] _exStage_WIRE_3_instr = 32'h00000000;
	wire [31:0] _exStage_WIRE_3_imm = 32'h00000000;
	wire [31:0] _exStage_WIRE_3_rs1Data = 32'h00000000;
	wire [31:0] _exStage_WIRE_3_rs2Data = 32'h00000000;
	wire [31:0] _exStage_WIRE_3_memAddr = 32'h00000000;
	wire [31:0] _exStage_WIRE_3_memWdata = 32'h00000000;
	wire [31:0] _exStage_WIRE_3_memRdata = 32'h00000000;
	wire [31:0] _exStage_WIRE_3_aluResult = 32'h00000000;
	wire [31:0] _exStage_WIRE_4_0_pc = 32'h00000000;
	wire [31:0] _exStage_WIRE_4_0_instr = 32'h00000000;
	wire [31:0] _exStage_WIRE_4_0_imm = 32'h00000000;
	wire [31:0] _exStage_WIRE_4_0_rs1Data = 32'h00000000;
	wire [31:0] _exStage_WIRE_4_0_rs2Data = 32'h00000000;
	wire [31:0] _exStage_WIRE_4_0_memAddr = 32'h00000000;
	wire [31:0] _exStage_WIRE_4_0_memWdata = 32'h00000000;
	wire [31:0] _exStage_WIRE_4_0_memRdata = 32'h00000000;
	wire [31:0] _exStage_WIRE_4_0_aluResult = 32'h00000000;
	wire [31:0] _exStage_WIRE_4_1_pc = 32'h00000000;
	wire [31:0] _exStage_WIRE_4_1_instr = 32'h00000000;
	wire [31:0] _exStage_WIRE_4_1_imm = 32'h00000000;
	wire [31:0] _exStage_WIRE_4_1_rs1Data = 32'h00000000;
	wire [31:0] _exStage_WIRE_4_1_rs2Data = 32'h00000000;
	wire [31:0] _exStage_WIRE_4_1_memAddr = 32'h00000000;
	wire [31:0] _exStage_WIRE_4_1_memWdata = 32'h00000000;
	wire [31:0] _exStage_WIRE_4_1_memRdata = 32'h00000000;
	wire [31:0] _exStage_WIRE_4_1_aluResult = 32'h00000000;
	wire [31:0] _exStage_WIRE_4_2_pc = 32'h00000000;
	wire [31:0] _exStage_WIRE_4_2_instr = 32'h00000000;
	wire [31:0] _exStage_WIRE_4_2_imm = 32'h00000000;
	wire [31:0] _exStage_WIRE_4_2_rs1Data = 32'h00000000;
	wire [31:0] _exStage_WIRE_4_2_rs2Data = 32'h00000000;
	wire [31:0] _exStage_WIRE_4_2_memAddr = 32'h00000000;
	wire [31:0] _exStage_WIRE_4_2_memWdata = 32'h00000000;
	wire [31:0] _exStage_WIRE_4_2_memRdata = 32'h00000000;
	wire [31:0] _exStage_WIRE_4_2_aluResult = 32'h00000000;
	wire [31:0] _exStage_WIRE_4_3_pc = 32'h00000000;
	wire [31:0] _exStage_WIRE_4_3_instr = 32'h00000000;
	wire [31:0] _exStage_WIRE_4_3_imm = 32'h00000000;
	wire [31:0] _exStage_WIRE_4_3_rs1Data = 32'h00000000;
	wire [31:0] _exStage_WIRE_4_3_rs2Data = 32'h00000000;
	wire [31:0] _exStage_WIRE_4_3_memAddr = 32'h00000000;
	wire [31:0] _exStage_WIRE_4_3_memWdata = 32'h00000000;
	wire [31:0] _exStage_WIRE_4_3_memRdata = 32'h00000000;
	wire [31:0] _exStage_WIRE_4_3_aluResult = 32'h00000000;
	wire [31:0] _memStage_WIRE_pc = 32'h00000000;
	wire [31:0] _memStage_WIRE_instr = 32'h00000000;
	wire [31:0] _memStage_WIRE_imm = 32'h00000000;
	wire [31:0] _memStage_WIRE_rs1Data = 32'h00000000;
	wire [31:0] _memStage_WIRE_rs2Data = 32'h00000000;
	wire [31:0] _memStage_WIRE_memAddr = 32'h00000000;
	wire [31:0] _memStage_WIRE_memWdata = 32'h00000000;
	wire [31:0] _memStage_WIRE_memRdata = 32'h00000000;
	wire [31:0] _memStage_WIRE_aluResult = 32'h00000000;
	wire [31:0] _memStage_WIRE_1_pc = 32'h00000000;
	wire [31:0] _memStage_WIRE_1_instr = 32'h00000000;
	wire [31:0] _memStage_WIRE_1_imm = 32'h00000000;
	wire [31:0] _memStage_WIRE_1_rs1Data = 32'h00000000;
	wire [31:0] _memStage_WIRE_1_rs2Data = 32'h00000000;
	wire [31:0] _memStage_WIRE_1_memAddr = 32'h00000000;
	wire [31:0] _memStage_WIRE_1_memWdata = 32'h00000000;
	wire [31:0] _memStage_WIRE_1_memRdata = 32'h00000000;
	wire [31:0] _memStage_WIRE_1_aluResult = 32'h00000000;
	wire [31:0] _memStage_WIRE_2_pc = 32'h00000000;
	wire [31:0] _memStage_WIRE_2_instr = 32'h00000000;
	wire [31:0] _memStage_WIRE_2_imm = 32'h00000000;
	wire [31:0] _memStage_WIRE_2_rs1Data = 32'h00000000;
	wire [31:0] _memStage_WIRE_2_rs2Data = 32'h00000000;
	wire [31:0] _memStage_WIRE_2_memAddr = 32'h00000000;
	wire [31:0] _memStage_WIRE_2_memWdata = 32'h00000000;
	wire [31:0] _memStage_WIRE_2_memRdata = 32'h00000000;
	wire [31:0] _memStage_WIRE_2_aluResult = 32'h00000000;
	wire [31:0] _memStage_WIRE_3_pc = 32'h00000000;
	wire [31:0] _memStage_WIRE_3_instr = 32'h00000000;
	wire [31:0] _memStage_WIRE_3_imm = 32'h00000000;
	wire [31:0] _memStage_WIRE_3_rs1Data = 32'h00000000;
	wire [31:0] _memStage_WIRE_3_rs2Data = 32'h00000000;
	wire [31:0] _memStage_WIRE_3_memAddr = 32'h00000000;
	wire [31:0] _memStage_WIRE_3_memWdata = 32'h00000000;
	wire [31:0] _memStage_WIRE_3_memRdata = 32'h00000000;
	wire [31:0] _memStage_WIRE_3_aluResult = 32'h00000000;
	wire [31:0] _memStage_WIRE_4_0_pc = 32'h00000000;
	wire [31:0] _memStage_WIRE_4_0_instr = 32'h00000000;
	wire [31:0] _memStage_WIRE_4_0_imm = 32'h00000000;
	wire [31:0] _memStage_WIRE_4_0_rs1Data = 32'h00000000;
	wire [31:0] _memStage_WIRE_4_0_rs2Data = 32'h00000000;
	wire [31:0] _memStage_WIRE_4_0_memAddr = 32'h00000000;
	wire [31:0] _memStage_WIRE_4_0_memWdata = 32'h00000000;
	wire [31:0] _memStage_WIRE_4_0_memRdata = 32'h00000000;
	wire [31:0] _memStage_WIRE_4_0_aluResult = 32'h00000000;
	wire [31:0] _memStage_WIRE_4_1_pc = 32'h00000000;
	wire [31:0] _memStage_WIRE_4_1_instr = 32'h00000000;
	wire [31:0] _memStage_WIRE_4_1_imm = 32'h00000000;
	wire [31:0] _memStage_WIRE_4_1_rs1Data = 32'h00000000;
	wire [31:0] _memStage_WIRE_4_1_rs2Data = 32'h00000000;
	wire [31:0] _memStage_WIRE_4_1_memAddr = 32'h00000000;
	wire [31:0] _memStage_WIRE_4_1_memWdata = 32'h00000000;
	wire [31:0] _memStage_WIRE_4_1_memRdata = 32'h00000000;
	wire [31:0] _memStage_WIRE_4_1_aluResult = 32'h00000000;
	wire [31:0] _memStage_WIRE_4_2_pc = 32'h00000000;
	wire [31:0] _memStage_WIRE_4_2_instr = 32'h00000000;
	wire [31:0] _memStage_WIRE_4_2_imm = 32'h00000000;
	wire [31:0] _memStage_WIRE_4_2_rs1Data = 32'h00000000;
	wire [31:0] _memStage_WIRE_4_2_rs2Data = 32'h00000000;
	wire [31:0] _memStage_WIRE_4_2_memAddr = 32'h00000000;
	wire [31:0] _memStage_WIRE_4_2_memWdata = 32'h00000000;
	wire [31:0] _memStage_WIRE_4_2_memRdata = 32'h00000000;
	wire [31:0] _memStage_WIRE_4_2_aluResult = 32'h00000000;
	wire [31:0] _memStage_WIRE_4_3_pc = 32'h00000000;
	wire [31:0] _memStage_WIRE_4_3_instr = 32'h00000000;
	wire [31:0] _memStage_WIRE_4_3_imm = 32'h00000000;
	wire [31:0] _memStage_WIRE_4_3_rs1Data = 32'h00000000;
	wire [31:0] _memStage_WIRE_4_3_rs2Data = 32'h00000000;
	wire [31:0] _memStage_WIRE_4_3_memAddr = 32'h00000000;
	wire [31:0] _memStage_WIRE_4_3_memWdata = 32'h00000000;
	wire [31:0] _memStage_WIRE_4_3_memRdata = 32'h00000000;
	wire [31:0] _memStage_WIRE_4_3_aluResult = 32'h00000000;
	wire [31:0] _ifWire_WIRE_pc = 32'h00000000;
	wire [31:0] _ifWire_WIRE_instr = 32'h00000000;
	wire [31:0] _ifWire_WIRE_imm = 32'h00000000;
	wire [31:0] _ifWire_WIRE_rs1Data = 32'h00000000;
	wire [31:0] _ifWire_WIRE_rs2Data = 32'h00000000;
	wire [31:0] _ifWire_WIRE_memAddr = 32'h00000000;
	wire [31:0] _ifWire_WIRE_memWdata = 32'h00000000;
	wire [31:0] _ifWire_WIRE_memRdata = 32'h00000000;
	wire [31:0] _ifWire_WIRE_aluResult = 32'h00000000;
	wire [31:0] ifWire_imm = 32'h00000000;
	wire [31:0] ifWire_rs1Data = 32'h00000000;
	wire [31:0] ifWire_rs2Data = 32'h00000000;
	wire [31:0] ifWire_memAddr = 32'h00000000;
	wire [31:0] ifWire_memWdata = 32'h00000000;
	wire [31:0] ifWire_memRdata = 32'h00000000;
	wire [31:0] ifWire_aluResult = 32'h00000000;
	wire [31:0] _decWire_WIRE_pc = 32'h00000000;
	wire [31:0] _decWire_WIRE_instr = 32'h00000000;
	wire [31:0] _decWire_WIRE_imm = 32'h00000000;
	wire [31:0] _decWire_WIRE_rs1Data = 32'h00000000;
	wire [31:0] _decWire_WIRE_rs2Data = 32'h00000000;
	wire [31:0] _decWire_WIRE_memAddr = 32'h00000000;
	wire [31:0] _decWire_WIRE_memWdata = 32'h00000000;
	wire [31:0] _decWire_WIRE_memRdata = 32'h00000000;
	wire [31:0] _decWire_WIRE_aluResult = 32'h00000000;
	wire [31:0] _exWire_WIRE_pc = 32'h00000000;
	wire [31:0] _exWire_WIRE_instr = 32'h00000000;
	wire [31:0] _exWire_WIRE_imm = 32'h00000000;
	wire [31:0] _exWire_WIRE_rs1Data = 32'h00000000;
	wire [31:0] _exWire_WIRE_rs2Data = 32'h00000000;
	wire [31:0] _exWire_WIRE_memAddr = 32'h00000000;
	wire [31:0] _exWire_WIRE_memWdata = 32'h00000000;
	wire [31:0] _exWire_WIRE_memRdata = 32'h00000000;
	wire [31:0] _exWire_WIRE_aluResult = 32'h00000000;
	wire [31:0] _memWire_WIRE_pc = 32'h00000000;
	wire [31:0] _memWire_WIRE_instr = 32'h00000000;
	wire [31:0] _memWire_WIRE_imm = 32'h00000000;
	wire [31:0] _memWire_WIRE_rs1Data = 32'h00000000;
	wire [31:0] _memWire_WIRE_rs2Data = 32'h00000000;
	wire [31:0] _memWire_WIRE_memAddr = 32'h00000000;
	wire [31:0] _memWire_WIRE_memWdata = 32'h00000000;
	wire [31:0] _memWire_WIRE_memRdata = 32'h00000000;
	wire [31:0] _memWire_WIRE_aluResult = 32'h00000000;
	wire [31:0] memWire_memAddr;
	wire [31:0] memWire_memWdata;
	wire [31:0] memWire_memRdata = io_memRdata_0;
	wire _io_memWe_T;
	reg [1:0] currentThread;
	wire [1:0] ifWire_threadId = currentThread;
	wire [2:0] _currentThread_T = {1'h0, currentThread} + 3'h1;
	wire [1:0] _currentThread_T_1 = _currentThread_T[1:0];
	reg [31:0] pcRegs_0;
	reg [31:0] pcRegs_1;
	reg [31:0] pcRegs_2;
	reg [31:0] pcRegs_3;
	reg [1:0] ifStage_0_threadId;
	reg ifStage_0_valid;
	reg [31:0] ifStage_0_pc;
	reg [31:0] ifStage_0_instr;
	reg [1:0] ifStage_1_threadId;
	reg ifStage_1_valid;
	reg [31:0] ifStage_1_pc;
	reg [31:0] ifStage_1_instr;
	reg [1:0] ifStage_2_threadId;
	reg ifStage_2_valid;
	reg [31:0] ifStage_2_pc;
	reg [31:0] ifStage_2_instr;
	reg [1:0] ifStage_3_threadId;
	reg ifStage_3_valid;
	reg [31:0] ifStage_3_pc;
	reg [31:0] ifStage_3_instr;
	reg [1:0] decStage_0_threadId;
	reg decStage_0_valid;
	reg [31:0] decStage_0_pc;
	reg [31:0] decStage_0_instr;
	reg decStage_0_isALU;
	reg decStage_0_isLoad;
	reg decStage_0_isStore;
	reg decStage_0_isBranch;
	reg decStage_0_isJAL;
	reg decStage_0_isJALR;
	reg decStage_0_isLUI;
	reg decStage_0_isAUIPC;
	reg decStage_0_isFence;
	reg decStage_0_isSystem;
	reg [4:0] decStage_0_aluOp;
	reg [31:0] decStage_0_imm;
	reg [4:0] decStage_0_rs1;
	reg [4:0] decStage_0_rs2;
	reg [4:0] decStage_0_rd;
	reg [31:0] decStage_0_rs1Data;
	reg [31:0] decStage_0_rs2Data;
	reg [31:0] decStage_0_memAddr;
	reg [31:0] decStage_0_memWdata;
	reg [31:0] decStage_0_memRdata;
	reg [31:0] decStage_0_aluResult;
	reg [1:0] decStage_1_threadId;
	reg decStage_1_valid;
	reg [31:0] decStage_1_pc;
	reg [31:0] decStage_1_instr;
	reg decStage_1_isALU;
	reg decStage_1_isLoad;
	reg decStage_1_isStore;
	reg decStage_1_isBranch;
	reg decStage_1_isJAL;
	reg decStage_1_isJALR;
	reg decStage_1_isLUI;
	reg decStage_1_isAUIPC;
	reg decStage_1_isFence;
	reg decStage_1_isSystem;
	reg [4:0] decStage_1_aluOp;
	reg [31:0] decStage_1_imm;
	reg [4:0] decStage_1_rs1;
	reg [4:0] decStage_1_rs2;
	reg [4:0] decStage_1_rd;
	reg [31:0] decStage_1_rs1Data;
	reg [31:0] decStage_1_rs2Data;
	reg [31:0] decStage_1_memAddr;
	reg [31:0] decStage_1_memWdata;
	reg [31:0] decStage_1_memRdata;
	reg [31:0] decStage_1_aluResult;
	reg [1:0] decStage_2_threadId;
	reg decStage_2_valid;
	reg [31:0] decStage_2_pc;
	reg [31:0] decStage_2_instr;
	reg decStage_2_isALU;
	reg decStage_2_isLoad;
	reg decStage_2_isStore;
	reg decStage_2_isBranch;
	reg decStage_2_isJAL;
	reg decStage_2_isJALR;
	reg decStage_2_isLUI;
	reg decStage_2_isAUIPC;
	reg decStage_2_isFence;
	reg decStage_2_isSystem;
	reg [4:0] decStage_2_aluOp;
	reg [31:0] decStage_2_imm;
	reg [4:0] decStage_2_rs1;
	reg [4:0] decStage_2_rs2;
	reg [4:0] decStage_2_rd;
	reg [31:0] decStage_2_rs1Data;
	reg [31:0] decStage_2_rs2Data;
	reg [31:0] decStage_2_memAddr;
	reg [31:0] decStage_2_memWdata;
	reg [31:0] decStage_2_memRdata;
	reg [31:0] decStage_2_aluResult;
	reg [1:0] decStage_3_threadId;
	reg decStage_3_valid;
	reg [31:0] decStage_3_pc;
	reg [31:0] decStage_3_instr;
	reg decStage_3_isALU;
	reg decStage_3_isLoad;
	reg decStage_3_isStore;
	reg decStage_3_isBranch;
	reg decStage_3_isJAL;
	reg decStage_3_isJALR;
	reg decStage_3_isLUI;
	reg decStage_3_isAUIPC;
	reg decStage_3_isFence;
	reg decStage_3_isSystem;
	reg [4:0] decStage_3_aluOp;
	reg [31:0] decStage_3_imm;
	reg [4:0] decStage_3_rs1;
	reg [4:0] decStage_3_rs2;
	reg [4:0] decStage_3_rd;
	reg [31:0] decStage_3_rs1Data;
	reg [31:0] decStage_3_rs2Data;
	reg [31:0] decStage_3_memAddr;
	reg [31:0] decStage_3_memWdata;
	reg [31:0] decStage_3_memRdata;
	reg [31:0] decStage_3_aluResult;
	reg [1:0] exStage_0_threadId;
	reg exStage_0_valid;
	reg [31:0] exStage_0_pc;
	reg [31:0] exStage_0_instr;
	reg exStage_0_isALU;
	reg exStage_0_isLoad;
	reg exStage_0_isStore;
	reg exStage_0_isBranch;
	reg exStage_0_isJAL;
	reg exStage_0_isJALR;
	reg exStage_0_isLUI;
	reg exStage_0_isAUIPC;
	reg exStage_0_isFence;
	reg exStage_0_isSystem;
	reg [4:0] exStage_0_aluOp;
	reg [31:0] exStage_0_imm;
	reg [4:0] exStage_0_rs1;
	reg [4:0] exStage_0_rs2;
	reg [4:0] exStage_0_rd;
	reg [31:0] exStage_0_rs1Data;
	reg [31:0] exStage_0_rs2Data;
	reg [31:0] exStage_0_memAddr;
	reg [31:0] exStage_0_memWdata;
	reg [31:0] exStage_0_memRdata;
	reg [31:0] exStage_0_aluResult;
	reg [1:0] exStage_1_threadId;
	reg exStage_1_valid;
	reg [31:0] exStage_1_pc;
	reg [31:0] exStage_1_instr;
	reg exStage_1_isALU;
	reg exStage_1_isLoad;
	reg exStage_1_isStore;
	reg exStage_1_isBranch;
	reg exStage_1_isJAL;
	reg exStage_1_isJALR;
	reg exStage_1_isLUI;
	reg exStage_1_isAUIPC;
	reg exStage_1_isFence;
	reg exStage_1_isSystem;
	reg [4:0] exStage_1_aluOp;
	reg [31:0] exStage_1_imm;
	reg [4:0] exStage_1_rs1;
	reg [4:0] exStage_1_rs2;
	reg [4:0] exStage_1_rd;
	reg [31:0] exStage_1_rs1Data;
	reg [31:0] exStage_1_rs2Data;
	reg [31:0] exStage_1_memAddr;
	reg [31:0] exStage_1_memWdata;
	reg [31:0] exStage_1_memRdata;
	reg [31:0] exStage_1_aluResult;
	reg [1:0] exStage_2_threadId;
	reg exStage_2_valid;
	reg [31:0] exStage_2_pc;
	reg [31:0] exStage_2_instr;
	reg exStage_2_isALU;
	reg exStage_2_isLoad;
	reg exStage_2_isStore;
	reg exStage_2_isBranch;
	reg exStage_2_isJAL;
	reg exStage_2_isJALR;
	reg exStage_2_isLUI;
	reg exStage_2_isAUIPC;
	reg exStage_2_isFence;
	reg exStage_2_isSystem;
	reg [4:0] exStage_2_aluOp;
	reg [31:0] exStage_2_imm;
	reg [4:0] exStage_2_rs1;
	reg [4:0] exStage_2_rs2;
	reg [4:0] exStage_2_rd;
	reg [31:0] exStage_2_rs1Data;
	reg [31:0] exStage_2_rs2Data;
	reg [31:0] exStage_2_memAddr;
	reg [31:0] exStage_2_memWdata;
	reg [31:0] exStage_2_memRdata;
	reg [31:0] exStage_2_aluResult;
	reg [1:0] exStage_3_threadId;
	reg exStage_3_valid;
	reg [31:0] exStage_3_pc;
	reg [31:0] exStage_3_instr;
	reg exStage_3_isALU;
	reg exStage_3_isLoad;
	reg exStage_3_isStore;
	reg exStage_3_isBranch;
	reg exStage_3_isJAL;
	reg exStage_3_isJALR;
	reg exStage_3_isLUI;
	reg exStage_3_isAUIPC;
	reg exStage_3_isFence;
	reg exStage_3_isSystem;
	reg [4:0] exStage_3_aluOp;
	reg [31:0] exStage_3_imm;
	reg [4:0] exStage_3_rs1;
	reg [4:0] exStage_3_rs2;
	reg [4:0] exStage_3_rd;
	reg [31:0] exStage_3_rs1Data;
	reg [31:0] exStage_3_rs2Data;
	reg [31:0] exStage_3_memAddr;
	reg [31:0] exStage_3_memWdata;
	reg [31:0] exStage_3_memRdata;
	reg [31:0] exStage_3_aluResult;
	reg [1:0] memStage_0_threadId;
	reg memStage_0_valid;
	reg [31:0] memStage_0_pc;
	reg [31:0] memStage_0_instr;
	reg memStage_0_isALU;
	reg memStage_0_isLoad;
	reg memStage_0_isStore;
	reg memStage_0_isBranch;
	reg memStage_0_isJAL;
	reg memStage_0_isJALR;
	reg memStage_0_isLUI;
	reg memStage_0_isAUIPC;
	reg memStage_0_isFence;
	reg memStage_0_isSystem;
	reg [4:0] memStage_0_aluOp;
	reg [31:0] memStage_0_imm;
	reg [4:0] memStage_0_rs1;
	reg [4:0] memStage_0_rs2;
	reg [4:0] memStage_0_rd;
	reg [31:0] memStage_0_rs1Data;
	reg [31:0] memStage_0_rs2Data;
	reg [31:0] memStage_0_memAddr;
	reg [31:0] memStage_0_memWdata;
	reg [31:0] memStage_0_memRdata;
	reg [31:0] memStage_0_aluResult;
	reg [1:0] memStage_1_threadId;
	reg memStage_1_valid;
	reg [31:0] memStage_1_pc;
	reg [31:0] memStage_1_instr;
	reg memStage_1_isALU;
	reg memStage_1_isLoad;
	reg memStage_1_isStore;
	reg memStage_1_isBranch;
	reg memStage_1_isJAL;
	reg memStage_1_isJALR;
	reg memStage_1_isLUI;
	reg memStage_1_isAUIPC;
	reg memStage_1_isFence;
	reg memStage_1_isSystem;
	reg [4:0] memStage_1_aluOp;
	reg [31:0] memStage_1_imm;
	reg [4:0] memStage_1_rs1;
	reg [4:0] memStage_1_rs2;
	reg [4:0] memStage_1_rd;
	reg [31:0] memStage_1_rs1Data;
	reg [31:0] memStage_1_rs2Data;
	reg [31:0] memStage_1_memAddr;
	reg [31:0] memStage_1_memWdata;
	reg [31:0] memStage_1_memRdata;
	reg [31:0] memStage_1_aluResult;
	reg [1:0] memStage_2_threadId;
	reg memStage_2_valid;
	reg [31:0] memStage_2_pc;
	reg [31:0] memStage_2_instr;
	reg memStage_2_isALU;
	reg memStage_2_isLoad;
	reg memStage_2_isStore;
	reg memStage_2_isBranch;
	reg memStage_2_isJAL;
	reg memStage_2_isJALR;
	reg memStage_2_isLUI;
	reg memStage_2_isAUIPC;
	reg memStage_2_isFence;
	reg memStage_2_isSystem;
	reg [4:0] memStage_2_aluOp;
	reg [31:0] memStage_2_imm;
	reg [4:0] memStage_2_rs1;
	reg [4:0] memStage_2_rs2;
	reg [4:0] memStage_2_rd;
	reg [31:0] memStage_2_rs1Data;
	reg [31:0] memStage_2_rs2Data;
	reg [31:0] memStage_2_memAddr;
	reg [31:0] memStage_2_memWdata;
	reg [31:0] memStage_2_memRdata;
	reg [31:0] memStage_2_aluResult;
	reg [1:0] memStage_3_threadId;
	reg memStage_3_valid;
	reg [31:0] memStage_3_pc;
	reg [31:0] memStage_3_instr;
	reg memStage_3_isALU;
	reg memStage_3_isLoad;
	reg memStage_3_isStore;
	reg memStage_3_isBranch;
	reg memStage_3_isJAL;
	reg memStage_3_isJALR;
	reg memStage_3_isLUI;
	reg memStage_3_isAUIPC;
	reg memStage_3_isFence;
	reg memStage_3_isSystem;
	reg [4:0] memStage_3_aluOp;
	reg [31:0] memStage_3_imm;
	reg [4:0] memStage_3_rs1;
	reg [4:0] memStage_3_rs2;
	reg [4:0] memStage_3_rd;
	reg [31:0] memStage_3_rs1Data;
	reg [31:0] memStage_3_rs2Data;
	reg [31:0] memStage_3_memAddr;
	reg [31:0] memStage_3_memWdata;
	reg [31:0] memStage_3_memRdata;
	reg [31:0] memStage_3_aluResult;
	wire [127:0] _GEN = {pcRegs_3, pcRegs_2, pcRegs_1, pcRegs_0};
	wire [31:0] ifWire_pc = _GEN[currentThread * 32+:32];
	wire [29:0] _ifWire_instr_T = ifWire_pc[31:2];
	wire [29:0] _ifWire_instr_WIRE = _ifWire_instr_T;
	wire [9:0] _ifWire_instr_T_1 = _ifWire_instr_WIRE[9:0];
	wire [32:0] _pcRegs_T = {1'h0, ifWire_pc} + 33'h000000004;
	wire [31:0] _pcRegs_T_1 = _pcRegs_T[31:0];
	wire [7:0] _GEN_0 = {decStage_3_threadId, decStage_2_threadId, decStage_1_threadId, decStage_0_threadId};
	wire [1:0] decWire_threadId = _GEN_0[currentThread * 2+:2];
	wire [3:0] _GEN_1 = {decStage_3_valid, decStage_2_valid, decStage_1_valid, decStage_0_valid};
	wire decWire_valid = _GEN_1[currentThread];
	wire [127:0] _GEN_2 = {decStage_3_pc, decStage_2_pc, decStage_1_pc, decStage_0_pc};
	wire [31:0] decWire_pc = _GEN_2[currentThread * 32+:32];
	wire [127:0] _GEN_3 = {decStage_3_instr, decStage_2_instr, decStage_1_instr, decStage_0_instr};
	wire [31:0] decWire_instr = _GEN_3[currentThread * 32+:32];
	wire [3:0] _GEN_4 = {decStage_3_isALU, decStage_2_isALU, decStage_1_isALU, decStage_0_isALU};
	wire [3:0] _GEN_5 = {decStage_3_isLoad, decStage_2_isLoad, decStage_1_isLoad, decStage_0_isLoad};
	wire [3:0] _GEN_6 = {decStage_3_isStore, decStage_2_isStore, decStage_1_isStore, decStage_0_isStore};
	wire [3:0] _GEN_7 = {decStage_3_isBranch, decStage_2_isBranch, decStage_1_isBranch, decStage_0_isBranch};
	wire decWire_isBranch = _GEN_7[currentThread];
	wire [3:0] _GEN_8 = {decStage_3_isJAL, decStage_2_isJAL, decStage_1_isJAL, decStage_0_isJAL};
	wire decWire_isJAL = _GEN_8[currentThread];
	wire [3:0] _GEN_9 = {decStage_3_isJALR, decStage_2_isJALR, decStage_1_isJALR, decStage_0_isJALR};
	wire decWire_isJALR = _GEN_9[currentThread];
	wire [3:0] _GEN_10 = {decStage_3_isLUI, decStage_2_isLUI, decStage_1_isLUI, decStage_0_isLUI};
	wire decWire_isLUI = _GEN_10[currentThread];
	wire [3:0] _GEN_11 = {decStage_3_isAUIPC, decStage_2_isAUIPC, decStage_1_isAUIPC, decStage_0_isAUIPC};
	wire decWire_isAUIPC = _GEN_11[currentThread];
	wire [3:0] _GEN_12 = {decStage_3_isFence, decStage_2_isFence, decStage_1_isFence, decStage_0_isFence};
	wire decWire_isFence = _GEN_12[currentThread];
	wire [3:0] _GEN_13 = {decStage_3_isSystem, decStage_2_isSystem, decStage_1_isSystem, decStage_0_isSystem};
	wire decWire_isSystem = _GEN_13[currentThread];
	wire [19:0] _GEN_14 = {decStage_3_aluOp, decStage_2_aluOp, decStage_1_aluOp, decStage_0_aluOp};
	wire [4:0] decWire_aluOp = _GEN_14[currentThread * 5+:5];
	wire [127:0] _GEN_15 = {decStage_3_imm, decStage_2_imm, decStage_1_imm, decStage_0_imm};
	wire [31:0] decWire_imm = _GEN_15[currentThread * 32+:32];
	wire [127:0] _GEN_16 = {decStage_3_memAddr, decStage_2_memAddr, decStage_1_memAddr, decStage_0_memAddr};
	wire [31:0] decWire_memAddr = _GEN_16[currentThread * 32+:32];
	wire [127:0] _GEN_17 = {decStage_3_memWdata, decStage_2_memWdata, decStage_1_memWdata, decStage_0_memWdata};
	wire [31:0] decWire_memWdata = _GEN_17[currentThread * 32+:32];
	wire [127:0] _GEN_18 = {decStage_3_memRdata, decStage_2_memRdata, decStage_1_memRdata, decStage_0_memRdata};
	wire [31:0] decWire_memRdata = _GEN_18[currentThread * 32+:32];
	wire [127:0] _GEN_19 = {decStage_3_aluResult, decStage_2_aluResult, decStage_1_aluResult, decStage_0_aluResult};
	wire [31:0] decWire_aluResult = _GEN_19[currentThread * 32+:32];
	wire [4:0] _decWire_rs1_T;
	wire [4:0] _decWire_rs2_T;
	wire [4:0] _decWire_rd_T;
	wire [6:0] opcode = decWire_instr[6:0];
	wire _T = opcode == 7'h33;
	wire decWire_isALU = _T | _GEN_4[currentThread];
	wire _T_1 = opcode == 7'h03;
	wire decWire_isLoad = (~_T & _T_1) | _GEN_5[currentThread];
	wire decWire_isStore = (~(_T | _T_1) & (opcode == 7'h23)) | _GEN_6[currentThread];
	assign _decWire_rs1_T = decWire_instr[19:15];
	wire [4:0] decWire_rs1 = _decWire_rs1_T;
	assign _decWire_rs2_T = decWire_instr[24:20];
	wire [4:0] decWire_rs2 = _decWire_rs2_T;
	assign _decWire_rd_T = decWire_instr[11:7];
	wire [4:0] decWire_rd = _decWire_rd_T;
	wire [7:0] _GEN_20 = {exStage_3_threadId, exStage_2_threadId, exStage_1_threadId, exStage_0_threadId};
	wire [1:0] exWire_threadId = _GEN_20[currentThread * 2+:2];
	wire [3:0] _GEN_21 = {exStage_3_valid, exStage_2_valid, exStage_1_valid, exStage_0_valid};
	wire exWire_valid = _GEN_21[currentThread];
	wire [127:0] _GEN_22 = {exStage_3_pc, exStage_2_pc, exStage_1_pc, exStage_0_pc};
	wire [31:0] exWire_pc = _GEN_22[currentThread * 32+:32];
	wire [127:0] _GEN_23 = {exStage_3_instr, exStage_2_instr, exStage_1_instr, exStage_0_instr};
	wire [31:0] exWire_instr = _GEN_23[currentThread * 32+:32];
	wire [3:0] _GEN_24 = {exStage_3_isALU, exStage_2_isALU, exStage_1_isALU, exStage_0_isALU};
	wire exWire_isALU = _GEN_24[currentThread];
	wire [3:0] _GEN_25 = {exStage_3_isLoad, exStage_2_isLoad, exStage_1_isLoad, exStage_0_isLoad};
	wire exWire_isLoad = _GEN_25[currentThread];
	wire [3:0] _GEN_26 = {exStage_3_isStore, exStage_2_isStore, exStage_1_isStore, exStage_0_isStore};
	wire exWire_isStore = _GEN_26[currentThread];
	wire [3:0] _GEN_27 = {exStage_3_isBranch, exStage_2_isBranch, exStage_1_isBranch, exStage_0_isBranch};
	wire exWire_isBranch = _GEN_27[currentThread];
	wire [3:0] _GEN_28 = {exStage_3_isJAL, exStage_2_isJAL, exStage_1_isJAL, exStage_0_isJAL};
	wire exWire_isJAL = _GEN_28[currentThread];
	wire [3:0] _GEN_29 = {exStage_3_isJALR, exStage_2_isJALR, exStage_1_isJALR, exStage_0_isJALR};
	wire exWire_isJALR = _GEN_29[currentThread];
	wire [3:0] _GEN_30 = {exStage_3_isLUI, exStage_2_isLUI, exStage_1_isLUI, exStage_0_isLUI};
	wire exWire_isLUI = _GEN_30[currentThread];
	wire [3:0] _GEN_31 = {exStage_3_isAUIPC, exStage_2_isAUIPC, exStage_1_isAUIPC, exStage_0_isAUIPC};
	wire exWire_isAUIPC = _GEN_31[currentThread];
	wire [3:0] _GEN_32 = {exStage_3_isFence, exStage_2_isFence, exStage_1_isFence, exStage_0_isFence};
	wire exWire_isFence = _GEN_32[currentThread];
	wire [3:0] _GEN_33 = {exStage_3_isSystem, exStage_2_isSystem, exStage_1_isSystem, exStage_0_isSystem};
	wire exWire_isSystem = _GEN_33[currentThread];
	wire [19:0] _GEN_34 = {exStage_3_aluOp, exStage_2_aluOp, exStage_1_aluOp, exStage_0_aluOp};
	wire [4:0] exWire_aluOp = _GEN_34[currentThread * 5+:5];
	wire [127:0] _GEN_35 = {exStage_3_imm, exStage_2_imm, exStage_1_imm, exStage_0_imm};
	wire [31:0] exWire_imm = _GEN_35[currentThread * 32+:32];
	wire [19:0] _GEN_36 = {exStage_3_rs1, exStage_2_rs1, exStage_1_rs1, exStage_0_rs1};
	wire [4:0] exWire_rs1 = _GEN_36[currentThread * 5+:5];
	wire [19:0] _GEN_37 = {exStage_3_rs2, exStage_2_rs2, exStage_1_rs2, exStage_0_rs2};
	wire [4:0] exWire_rs2 = _GEN_37[currentThread * 5+:5];
	wire [19:0] _GEN_38 = {exStage_3_rd, exStage_2_rd, exStage_1_rd, exStage_0_rd};
	wire [4:0] exWire_rd = _GEN_38[currentThread * 5+:5];
	wire [127:0] _GEN_39 = {exStage_3_rs1Data, exStage_2_rs1Data, exStage_1_rs1Data, exStage_0_rs1Data};
	wire [31:0] exWire_rs1Data = _GEN_39[currentThread * 32+:32];
	wire [127:0] _GEN_40 = {exStage_3_rs2Data, exStage_2_rs2Data, exStage_1_rs2Data, exStage_0_rs2Data};
	wire [31:0] exWire_rs2Data = _GEN_40[currentThread * 32+:32];
	wire [127:0] _GEN_41 = {exStage_3_memAddr, exStage_2_memAddr, exStage_1_memAddr, exStage_0_memAddr};
	wire [127:0] _GEN_42 = {exStage_3_memWdata, exStage_2_memWdata, exStage_1_memWdata, exStage_0_memWdata};
	wire [127:0] _GEN_43 = {exStage_3_memRdata, exStage_2_memRdata, exStage_1_memRdata, exStage_0_memRdata};
	wire [31:0] exWire_memRdata = _GEN_43[currentThread * 32+:32];
	wire _T_3 = exWire_isLoad | exWire_isStore;
	wire [32:0] _exWire_memAddr_T = {1'h0, exWire_rs1Data} + {1'h0, exWire_imm};
	wire [31:0] _exWire_memAddr_T_1 = _exWire_memAddr_T[31:0];
	wire [31:0] exWire_memAddr = (_T_3 ? _exWire_memAddr_T_1 : _GEN_41[currentThread * 32+:32]);
	wire [31:0] exWire_memWdata = (_T_3 ? exWire_rs2Data : _GEN_42[currentThread * 32+:32]);
	wire [7:0] _GEN_44 = {memStage_3_threadId, memStage_2_threadId, memStage_1_threadId, memStage_0_threadId};
	wire [1:0] memWire_threadId = _GEN_44[currentThread * 2+:2];
	wire [3:0] _GEN_45 = {memStage_3_valid, memStage_2_valid, memStage_1_valid, memStage_0_valid};
	wire memWire_valid = _GEN_45[currentThread];
	wire [127:0] _GEN_46 = {memStage_3_pc, memStage_2_pc, memStage_1_pc, memStage_0_pc};
	wire [31:0] memWire_pc = _GEN_46[currentThread * 32+:32];
	wire [127:0] _GEN_47 = {memStage_3_instr, memStage_2_instr, memStage_1_instr, memStage_0_instr};
	wire [31:0] memWire_instr = _GEN_47[currentThread * 32+:32];
	wire [3:0] _GEN_48 = {memStage_3_isALU, memStage_2_isALU, memStage_1_isALU, memStage_0_isALU};
	wire memWire_isALU = _GEN_48[currentThread];
	wire [3:0] _GEN_49 = {memStage_3_isLoad, memStage_2_isLoad, memStage_1_isLoad, memStage_0_isLoad};
	wire memWire_isLoad = _GEN_49[currentThread];
	wire [3:0] _GEN_50 = {memStage_3_isStore, memStage_2_isStore, memStage_1_isStore, memStage_0_isStore};
	wire memWire_isStore = _GEN_50[currentThread];
	wire [3:0] _GEN_51 = {memStage_3_isBranch, memStage_2_isBranch, memStage_1_isBranch, memStage_0_isBranch};
	wire memWire_isBranch = _GEN_51[currentThread];
	wire [3:0] _GEN_52 = {memStage_3_isJAL, memStage_2_isJAL, memStage_1_isJAL, memStage_0_isJAL};
	wire memWire_isJAL = _GEN_52[currentThread];
	wire [3:0] _GEN_53 = {memStage_3_isJALR, memStage_2_isJALR, memStage_1_isJALR, memStage_0_isJALR};
	wire memWire_isJALR = _GEN_53[currentThread];
	wire [3:0] _GEN_54 = {memStage_3_isLUI, memStage_2_isLUI, memStage_1_isLUI, memStage_0_isLUI};
	wire memWire_isLUI = _GEN_54[currentThread];
	wire [3:0] _GEN_55 = {memStage_3_isAUIPC, memStage_2_isAUIPC, memStage_1_isAUIPC, memStage_0_isAUIPC};
	wire memWire_isAUIPC = _GEN_55[currentThread];
	wire [3:0] _GEN_56 = {memStage_3_isFence, memStage_2_isFence, memStage_1_isFence, memStage_0_isFence};
	wire memWire_isFence = _GEN_56[currentThread];
	wire [3:0] _GEN_57 = {memStage_3_isSystem, memStage_2_isSystem, memStage_1_isSystem, memStage_0_isSystem};
	wire memWire_isSystem = _GEN_57[currentThread];
	wire [19:0] _GEN_58 = {memStage_3_aluOp, memStage_2_aluOp, memStage_1_aluOp, memStage_0_aluOp};
	wire [4:0] memWire_aluOp = _GEN_58[currentThread * 5+:5];
	wire [127:0] _GEN_59 = {memStage_3_imm, memStage_2_imm, memStage_1_imm, memStage_0_imm};
	wire [31:0] memWire_imm = _GEN_59[currentThread * 32+:32];
	wire [19:0] _GEN_60 = {memStage_3_rs1, memStage_2_rs1, memStage_1_rs1, memStage_0_rs1};
	wire [4:0] memWire_rs1 = _GEN_60[currentThread * 5+:5];
	wire [19:0] _GEN_61 = {memStage_3_rs2, memStage_2_rs2, memStage_1_rs2, memStage_0_rs2};
	wire [4:0] memWire_rs2 = _GEN_61[currentThread * 5+:5];
	wire [19:0] _GEN_62 = {memStage_3_rd, memStage_2_rd, memStage_1_rd, memStage_0_rd};
	wire [4:0] memWire_rd = _GEN_62[currentThread * 5+:5];
	wire [127:0] _GEN_63 = {memStage_3_rs1Data, memStage_2_rs1Data, memStage_1_rs1Data, memStage_0_rs1Data};
	wire [31:0] memWire_rs1Data = _GEN_63[currentThread * 32+:32];
	wire [127:0] _GEN_64 = {memStage_3_rs2Data, memStage_2_rs2Data, memStage_1_rs2Data, memStage_0_rs2Data};
	wire [31:0] memWire_rs2Data = _GEN_64[currentThread * 32+:32];
	wire [127:0] _GEN_65 = {memStage_3_memAddr, memStage_2_memAddr, memStage_1_memAddr, memStage_0_memAddr};
	assign memWire_memAddr = _GEN_65[currentThread * 32+:32];
	wire [127:0] _GEN_66 = {memStage_3_memWdata, memStage_2_memWdata, memStage_1_memWdata, memStage_0_memWdata};
	assign memWire_memWdata = _GEN_66[currentThread * 32+:32];
	wire [127:0] _GEN_67 = {memStage_3_aluResult, memStage_2_aluResult, memStage_1_aluResult, memStage_0_aluResult};
	wire [31:0] memWire_aluResult = _GEN_67[currentThread * 32+:32];
	wire [31:0] io_memAddr_0 = memWire_memAddr;
	wire [31:0] io_memWdata_0 = memWire_memWdata;
	assign _io_memWe_T = memWire_isStore & memWire_valid;
	wire io_memWe_0 = _io_memWe_T;
	wire [31:0] wbData = (memWire_isLoad ? memWire_memRdata : memWire_aluResult);
	wire _regFile_io_wen_T = |memWire_rd;
	wire _regFile_io_wen_T_1 = memWire_valid & _regFile_io_wen_T;
	wire _regFile_io_wen_T_2 = memWire_isLoad | memWire_isALU;
	wire _regFile_io_wen_T_3 = _regFile_io_wen_T_1 & _regFile_io_wen_T_2;
	wire [31:0] ifWire_instr;
	wire [31:0] decWire_rs1Data;
	wire [31:0] decWire_rs2Data;
	wire [31:0] exWire_aluResult;
	always @(posedge clock)
		if (reset) begin
			currentThread <= 2'h0;
			pcRegs_0 <= 32'h00000000;
			pcRegs_1 <= 32'h00000000;
			pcRegs_2 <= 32'h00000000;
			pcRegs_3 <= 32'h00000000;
			ifStage_0_threadId <= 2'h0;
			ifStage_0_valid <= 1'h0;
			ifStage_0_pc <= 32'h00000000;
			ifStage_0_instr <= 32'h00000000;
			ifStage_1_threadId <= 2'h0;
			ifStage_1_valid <= 1'h0;
			ifStage_1_pc <= 32'h00000000;
			ifStage_1_instr <= 32'h00000000;
			ifStage_2_threadId <= 2'h0;
			ifStage_2_valid <= 1'h0;
			ifStage_2_pc <= 32'h00000000;
			ifStage_2_instr <= 32'h00000000;
			ifStage_3_threadId <= 2'h0;
			ifStage_3_valid <= 1'h0;
			ifStage_3_pc <= 32'h00000000;
			ifStage_3_instr <= 32'h00000000;
			decStage_0_threadId <= 2'h0;
			decStage_0_valid <= 1'h0;
			decStage_0_pc <= 32'h00000000;
			decStage_0_instr <= 32'h00000000;
			decStage_0_isALU <= 1'h0;
			decStage_0_isLoad <= 1'h0;
			decStage_0_isStore <= 1'h0;
			decStage_0_isBranch <= 1'h0;
			decStage_0_isJAL <= 1'h0;
			decStage_0_isJALR <= 1'h0;
			decStage_0_isLUI <= 1'h0;
			decStage_0_isAUIPC <= 1'h0;
			decStage_0_isFence <= 1'h0;
			decStage_0_isSystem <= 1'h0;
			decStage_0_aluOp <= 5'h00;
			decStage_0_imm <= 32'h00000000;
			decStage_0_rs1 <= 5'h00;
			decStage_0_rs2 <= 5'h00;
			decStage_0_rd <= 5'h00;
			decStage_0_rs1Data <= 32'h00000000;
			decStage_0_rs2Data <= 32'h00000000;
			decStage_0_memAddr <= 32'h00000000;
			decStage_0_memWdata <= 32'h00000000;
			decStage_0_memRdata <= 32'h00000000;
			decStage_0_aluResult <= 32'h00000000;
			decStage_1_threadId <= 2'h0;
			decStage_1_valid <= 1'h0;
			decStage_1_pc <= 32'h00000000;
			decStage_1_instr <= 32'h00000000;
			decStage_1_isALU <= 1'h0;
			decStage_1_isLoad <= 1'h0;
			decStage_1_isStore <= 1'h0;
			decStage_1_isBranch <= 1'h0;
			decStage_1_isJAL <= 1'h0;
			decStage_1_isJALR <= 1'h0;
			decStage_1_isLUI <= 1'h0;
			decStage_1_isAUIPC <= 1'h0;
			decStage_1_isFence <= 1'h0;
			decStage_1_isSystem <= 1'h0;
			decStage_1_aluOp <= 5'h00;
			decStage_1_imm <= 32'h00000000;
			decStage_1_rs1 <= 5'h00;
			decStage_1_rs2 <= 5'h00;
			decStage_1_rd <= 5'h00;
			decStage_1_rs1Data <= 32'h00000000;
			decStage_1_rs2Data <= 32'h00000000;
			decStage_1_memAddr <= 32'h00000000;
			decStage_1_memWdata <= 32'h00000000;
			decStage_1_memRdata <= 32'h00000000;
			decStage_1_aluResult <= 32'h00000000;
			decStage_2_threadId <= 2'h0;
			decStage_2_valid <= 1'h0;
			decStage_2_pc <= 32'h00000000;
			decStage_2_instr <= 32'h00000000;
			decStage_2_isALU <= 1'h0;
			decStage_2_isLoad <= 1'h0;
			decStage_2_isStore <= 1'h0;
			decStage_2_isBranch <= 1'h0;
			decStage_2_isJAL <= 1'h0;
			decStage_2_isJALR <= 1'h0;
			decStage_2_isLUI <= 1'h0;
			decStage_2_isAUIPC <= 1'h0;
			decStage_2_isFence <= 1'h0;
			decStage_2_isSystem <= 1'h0;
			decStage_2_aluOp <= 5'h00;
			decStage_2_imm <= 32'h00000000;
			decStage_2_rs1 <= 5'h00;
			decStage_2_rs2 <= 5'h00;
			decStage_2_rd <= 5'h00;
			decStage_2_rs1Data <= 32'h00000000;
			decStage_2_rs2Data <= 32'h00000000;
			decStage_2_memAddr <= 32'h00000000;
			decStage_2_memWdata <= 32'h00000000;
			decStage_2_memRdata <= 32'h00000000;
			decStage_2_aluResult <= 32'h00000000;
			decStage_3_threadId <= 2'h0;
			decStage_3_valid <= 1'h0;
			decStage_3_pc <= 32'h00000000;
			decStage_3_instr <= 32'h00000000;
			decStage_3_isALU <= 1'h0;
			decStage_3_isLoad <= 1'h0;
			decStage_3_isStore <= 1'h0;
			decStage_3_isBranch <= 1'h0;
			decStage_3_isJAL <= 1'h0;
			decStage_3_isJALR <= 1'h0;
			decStage_3_isLUI <= 1'h0;
			decStage_3_isAUIPC <= 1'h0;
			decStage_3_isFence <= 1'h0;
			decStage_3_isSystem <= 1'h0;
			decStage_3_aluOp <= 5'h00;
			decStage_3_imm <= 32'h00000000;
			decStage_3_rs1 <= 5'h00;
			decStage_3_rs2 <= 5'h00;
			decStage_3_rd <= 5'h00;
			decStage_3_rs1Data <= 32'h00000000;
			decStage_3_rs2Data <= 32'h00000000;
			decStage_3_memAddr <= 32'h00000000;
			decStage_3_memWdata <= 32'h00000000;
			decStage_3_memRdata <= 32'h00000000;
			decStage_3_aluResult <= 32'h00000000;
			exStage_0_threadId <= 2'h0;
			exStage_0_valid <= 1'h0;
			exStage_0_pc <= 32'h00000000;
			exStage_0_instr <= 32'h00000000;
			exStage_0_isALU <= 1'h0;
			exStage_0_isLoad <= 1'h0;
			exStage_0_isStore <= 1'h0;
			exStage_0_isBranch <= 1'h0;
			exStage_0_isJAL <= 1'h0;
			exStage_0_isJALR <= 1'h0;
			exStage_0_isLUI <= 1'h0;
			exStage_0_isAUIPC <= 1'h0;
			exStage_0_isFence <= 1'h0;
			exStage_0_isSystem <= 1'h0;
			exStage_0_aluOp <= 5'h00;
			exStage_0_imm <= 32'h00000000;
			exStage_0_rs1 <= 5'h00;
			exStage_0_rs2 <= 5'h00;
			exStage_0_rd <= 5'h00;
			exStage_0_rs1Data <= 32'h00000000;
			exStage_0_rs2Data <= 32'h00000000;
			exStage_0_memAddr <= 32'h00000000;
			exStage_0_memWdata <= 32'h00000000;
			exStage_0_memRdata <= 32'h00000000;
			exStage_0_aluResult <= 32'h00000000;
			exStage_1_threadId <= 2'h0;
			exStage_1_valid <= 1'h0;
			exStage_1_pc <= 32'h00000000;
			exStage_1_instr <= 32'h00000000;
			exStage_1_isALU <= 1'h0;
			exStage_1_isLoad <= 1'h0;
			exStage_1_isStore <= 1'h0;
			exStage_1_isBranch <= 1'h0;
			exStage_1_isJAL <= 1'h0;
			exStage_1_isJALR <= 1'h0;
			exStage_1_isLUI <= 1'h0;
			exStage_1_isAUIPC <= 1'h0;
			exStage_1_isFence <= 1'h0;
			exStage_1_isSystem <= 1'h0;
			exStage_1_aluOp <= 5'h00;
			exStage_1_imm <= 32'h00000000;
			exStage_1_rs1 <= 5'h00;
			exStage_1_rs2 <= 5'h00;
			exStage_1_rd <= 5'h00;
			exStage_1_rs1Data <= 32'h00000000;
			exStage_1_rs2Data <= 32'h00000000;
			exStage_1_memAddr <= 32'h00000000;
			exStage_1_memWdata <= 32'h00000000;
			exStage_1_memRdata <= 32'h00000000;
			exStage_1_aluResult <= 32'h00000000;
			exStage_2_threadId <= 2'h0;
			exStage_2_valid <= 1'h0;
			exStage_2_pc <= 32'h00000000;
			exStage_2_instr <= 32'h00000000;
			exStage_2_isALU <= 1'h0;
			exStage_2_isLoad <= 1'h0;
			exStage_2_isStore <= 1'h0;
			exStage_2_isBranch <= 1'h0;
			exStage_2_isJAL <= 1'h0;
			exStage_2_isJALR <= 1'h0;
			exStage_2_isLUI <= 1'h0;
			exStage_2_isAUIPC <= 1'h0;
			exStage_2_isFence <= 1'h0;
			exStage_2_isSystem <= 1'h0;
			exStage_2_aluOp <= 5'h00;
			exStage_2_imm <= 32'h00000000;
			exStage_2_rs1 <= 5'h00;
			exStage_2_rs2 <= 5'h00;
			exStage_2_rd <= 5'h00;
			exStage_2_rs1Data <= 32'h00000000;
			exStage_2_rs2Data <= 32'h00000000;
			exStage_2_memAddr <= 32'h00000000;
			exStage_2_memWdata <= 32'h00000000;
			exStage_2_memRdata <= 32'h00000000;
			exStage_2_aluResult <= 32'h00000000;
			exStage_3_threadId <= 2'h0;
			exStage_3_valid <= 1'h0;
			exStage_3_pc <= 32'h00000000;
			exStage_3_instr <= 32'h00000000;
			exStage_3_isALU <= 1'h0;
			exStage_3_isLoad <= 1'h0;
			exStage_3_isStore <= 1'h0;
			exStage_3_isBranch <= 1'h0;
			exStage_3_isJAL <= 1'h0;
			exStage_3_isJALR <= 1'h0;
			exStage_3_isLUI <= 1'h0;
			exStage_3_isAUIPC <= 1'h0;
			exStage_3_isFence <= 1'h0;
			exStage_3_isSystem <= 1'h0;
			exStage_3_aluOp <= 5'h00;
			exStage_3_imm <= 32'h00000000;
			exStage_3_rs1 <= 5'h00;
			exStage_3_rs2 <= 5'h00;
			exStage_3_rd <= 5'h00;
			exStage_3_rs1Data <= 32'h00000000;
			exStage_3_rs2Data <= 32'h00000000;
			exStage_3_memAddr <= 32'h00000000;
			exStage_3_memWdata <= 32'h00000000;
			exStage_3_memRdata <= 32'h00000000;
			exStage_3_aluResult <= 32'h00000000;
			memStage_0_threadId <= 2'h0;
			memStage_0_valid <= 1'h0;
			memStage_0_pc <= 32'h00000000;
			memStage_0_instr <= 32'h00000000;
			memStage_0_isALU <= 1'h0;
			memStage_0_isLoad <= 1'h0;
			memStage_0_isStore <= 1'h0;
			memStage_0_isBranch <= 1'h0;
			memStage_0_isJAL <= 1'h0;
			memStage_0_isJALR <= 1'h0;
			memStage_0_isLUI <= 1'h0;
			memStage_0_isAUIPC <= 1'h0;
			memStage_0_isFence <= 1'h0;
			memStage_0_isSystem <= 1'h0;
			memStage_0_aluOp <= 5'h00;
			memStage_0_imm <= 32'h00000000;
			memStage_0_rs1 <= 5'h00;
			memStage_0_rs2 <= 5'h00;
			memStage_0_rd <= 5'h00;
			memStage_0_rs1Data <= 32'h00000000;
			memStage_0_rs2Data <= 32'h00000000;
			memStage_0_memAddr <= 32'h00000000;
			memStage_0_memWdata <= 32'h00000000;
			memStage_0_memRdata <= 32'h00000000;
			memStage_0_aluResult <= 32'h00000000;
			memStage_1_threadId <= 2'h0;
			memStage_1_valid <= 1'h0;
			memStage_1_pc <= 32'h00000000;
			memStage_1_instr <= 32'h00000000;
			memStage_1_isALU <= 1'h0;
			memStage_1_isLoad <= 1'h0;
			memStage_1_isStore <= 1'h0;
			memStage_1_isBranch <= 1'h0;
			memStage_1_isJAL <= 1'h0;
			memStage_1_isJALR <= 1'h0;
			memStage_1_isLUI <= 1'h0;
			memStage_1_isAUIPC <= 1'h0;
			memStage_1_isFence <= 1'h0;
			memStage_1_isSystem <= 1'h0;
			memStage_1_aluOp <= 5'h00;
			memStage_1_imm <= 32'h00000000;
			memStage_1_rs1 <= 5'h00;
			memStage_1_rs2 <= 5'h00;
			memStage_1_rd <= 5'h00;
			memStage_1_rs1Data <= 32'h00000000;
			memStage_1_rs2Data <= 32'h00000000;
			memStage_1_memAddr <= 32'h00000000;
			memStage_1_memWdata <= 32'h00000000;
			memStage_1_memRdata <= 32'h00000000;
			memStage_1_aluResult <= 32'h00000000;
			memStage_2_threadId <= 2'h0;
			memStage_2_valid <= 1'h0;
			memStage_2_pc <= 32'h00000000;
			memStage_2_instr <= 32'h00000000;
			memStage_2_isALU <= 1'h0;
			memStage_2_isLoad <= 1'h0;
			memStage_2_isStore <= 1'h0;
			memStage_2_isBranch <= 1'h0;
			memStage_2_isJAL <= 1'h0;
			memStage_2_isJALR <= 1'h0;
			memStage_2_isLUI <= 1'h0;
			memStage_2_isAUIPC <= 1'h0;
			memStage_2_isFence <= 1'h0;
			memStage_2_isSystem <= 1'h0;
			memStage_2_aluOp <= 5'h00;
			memStage_2_imm <= 32'h00000000;
			memStage_2_rs1 <= 5'h00;
			memStage_2_rs2 <= 5'h00;
			memStage_2_rd <= 5'h00;
			memStage_2_rs1Data <= 32'h00000000;
			memStage_2_rs2Data <= 32'h00000000;
			memStage_2_memAddr <= 32'h00000000;
			memStage_2_memWdata <= 32'h00000000;
			memStage_2_memRdata <= 32'h00000000;
			memStage_2_aluResult <= 32'h00000000;
			memStage_3_threadId <= 2'h0;
			memStage_3_valid <= 1'h0;
			memStage_3_pc <= 32'h00000000;
			memStage_3_instr <= 32'h00000000;
			memStage_3_isALU <= 1'h0;
			memStage_3_isLoad <= 1'h0;
			memStage_3_isStore <= 1'h0;
			memStage_3_isBranch <= 1'h0;
			memStage_3_isJAL <= 1'h0;
			memStage_3_isJALR <= 1'h0;
			memStage_3_isLUI <= 1'h0;
			memStage_3_isAUIPC <= 1'h0;
			memStage_3_isFence <= 1'h0;
			memStage_3_isSystem <= 1'h0;
			memStage_3_aluOp <= 5'h00;
			memStage_3_imm <= 32'h00000000;
			memStage_3_rs1 <= 5'h00;
			memStage_3_rs2 <= 5'h00;
			memStage_3_rd <= 5'h00;
			memStage_3_rs1Data <= 32'h00000000;
			memStage_3_rs2Data <= 32'h00000000;
			memStage_3_memAddr <= 32'h00000000;
			memStage_3_memWdata <= 32'h00000000;
			memStage_3_memRdata <= 32'h00000000;
			memStage_3_aluResult <= 32'h00000000;
		end
		else begin : sv2v_autoblock_1
			reg _GEN_68;
			reg _GEN_69;
			reg _GEN_70;
			_GEN_68 = currentThread == 2'h0;
			_GEN_69 = currentThread == 2'h1;
			_GEN_70 = currentThread == 2'h2;
			currentThread <= _currentThread_T_1;
			if (_GEN_68) begin
				pcRegs_0 <= _pcRegs_T_1;
				ifStage_0_threadId <= ifWire_threadId;
				ifStage_0_pc <= ifWire_pc;
				ifStage_0_instr <= ifWire_instr;
				decStage_0_threadId <= decWire_threadId;
				decStage_0_valid <= decWire_valid;
				decStage_0_pc <= decWire_pc;
				decStage_0_instr <= decWire_instr;
				decStage_0_aluOp <= decWire_aluOp;
				decStage_0_imm <= decWire_imm;
				decStage_0_rs1 <= decWire_rs1;
				decStage_0_rs2 <= decWire_rs2;
				decStage_0_rd <= decWire_rd;
				decStage_0_rs1Data <= decWire_rs1Data;
				decStage_0_rs2Data <= decWire_rs2Data;
				decStage_0_memAddr <= decWire_memAddr;
				decStage_0_memWdata <= decWire_memWdata;
				decStage_0_memRdata <= decWire_memRdata;
				decStage_0_aluResult <= decWire_aluResult;
				exStage_0_threadId <= exWire_threadId;
				exStage_0_valid <= exWire_valid;
				exStage_0_pc <= exWire_pc;
				exStage_0_instr <= exWire_instr;
				exStage_0_isALU <= exWire_isALU;
				exStage_0_isLoad <= exWire_isLoad;
				exStage_0_isStore <= exWire_isStore;
				exStage_0_isBranch <= exWire_isBranch;
				exStage_0_isJAL <= exWire_isJAL;
				exStage_0_isJALR <= exWire_isJALR;
				exStage_0_isLUI <= exWire_isLUI;
				exStage_0_isAUIPC <= exWire_isAUIPC;
				exStage_0_isFence <= exWire_isFence;
				exStage_0_isSystem <= exWire_isSystem;
				exStage_0_aluOp <= exWire_aluOp;
				exStage_0_imm <= exWire_imm;
				exStage_0_rs1 <= exWire_rs1;
				exStage_0_rs2 <= exWire_rs2;
				exStage_0_rd <= exWire_rd;
				exStage_0_rs1Data <= exWire_rs1Data;
				exStage_0_rs2Data <= exWire_rs2Data;
				exStage_0_memAddr <= exWire_memAddr;
				exStage_0_memWdata <= exWire_memWdata;
				exStage_0_memRdata <= exWire_memRdata;
				exStage_0_aluResult <= exWire_aluResult;
				memStage_0_threadId <= memWire_threadId;
				memStage_0_valid <= memWire_valid;
				memStage_0_pc <= memWire_pc;
				memStage_0_instr <= memWire_instr;
				memStage_0_isALU <= memWire_isALU;
				memStage_0_isLoad <= memWire_isLoad;
				memStage_0_isStore <= memWire_isStore;
				memStage_0_isBranch <= memWire_isBranch;
				memStage_0_isJAL <= memWire_isJAL;
				memStage_0_isJALR <= memWire_isJALR;
				memStage_0_isLUI <= memWire_isLUI;
				memStage_0_isAUIPC <= memWire_isAUIPC;
				memStage_0_isFence <= memWire_isFence;
				memStage_0_isSystem <= memWire_isSystem;
				memStage_0_aluOp <= memWire_aluOp;
				memStage_0_imm <= memWire_imm;
				memStage_0_rs1 <= memWire_rs1;
				memStage_0_rs2 <= memWire_rs2;
				memStage_0_rd <= memWire_rd;
				memStage_0_rs1Data <= memWire_rs1Data;
				memStage_0_rs2Data <= memWire_rs2Data;
				memStage_0_memAddr <= memWire_memAddr;
				memStage_0_memWdata <= memWire_memWdata;
				memStage_0_memRdata <= memWire_memRdata;
				memStage_0_aluResult <= memWire_aluResult;
			end
			if (_GEN_69) begin
				pcRegs_1 <= _pcRegs_T_1;
				ifStage_1_threadId <= ifWire_threadId;
				ifStage_1_pc <= ifWire_pc;
				ifStage_1_instr <= ifWire_instr;
				decStage_1_threadId <= decWire_threadId;
				decStage_1_valid <= decWire_valid;
				decStage_1_pc <= decWire_pc;
				decStage_1_instr <= decWire_instr;
				decStage_1_aluOp <= decWire_aluOp;
				decStage_1_imm <= decWire_imm;
				decStage_1_rs1 <= decWire_rs1;
				decStage_1_rs2 <= decWire_rs2;
				decStage_1_rd <= decWire_rd;
				decStage_1_rs1Data <= decWire_rs1Data;
				decStage_1_rs2Data <= decWire_rs2Data;
				decStage_1_memAddr <= decWire_memAddr;
				decStage_1_memWdata <= decWire_memWdata;
				decStage_1_memRdata <= decWire_memRdata;
				decStage_1_aluResult <= decWire_aluResult;
				exStage_1_threadId <= exWire_threadId;
				exStage_1_valid <= exWire_valid;
				exStage_1_pc <= exWire_pc;
				exStage_1_instr <= exWire_instr;
				exStage_1_isALU <= exWire_isALU;
				exStage_1_isLoad <= exWire_isLoad;
				exStage_1_isStore <= exWire_isStore;
				exStage_1_isBranch <= exWire_isBranch;
				exStage_1_isJAL <= exWire_isJAL;
				exStage_1_isJALR <= exWire_isJALR;
				exStage_1_isLUI <= exWire_isLUI;
				exStage_1_isAUIPC <= exWire_isAUIPC;
				exStage_1_isFence <= exWire_isFence;
				exStage_1_isSystem <= exWire_isSystem;
				exStage_1_aluOp <= exWire_aluOp;
				exStage_1_imm <= exWire_imm;
				exStage_1_rs1 <= exWire_rs1;
				exStage_1_rs2 <= exWire_rs2;
				exStage_1_rd <= exWire_rd;
				exStage_1_rs1Data <= exWire_rs1Data;
				exStage_1_rs2Data <= exWire_rs2Data;
				exStage_1_memAddr <= exWire_memAddr;
				exStage_1_memWdata <= exWire_memWdata;
				exStage_1_memRdata <= exWire_memRdata;
				exStage_1_aluResult <= exWire_aluResult;
				memStage_1_threadId <= memWire_threadId;
				memStage_1_valid <= memWire_valid;
				memStage_1_pc <= memWire_pc;
				memStage_1_instr <= memWire_instr;
				memStage_1_isALU <= memWire_isALU;
				memStage_1_isLoad <= memWire_isLoad;
				memStage_1_isStore <= memWire_isStore;
				memStage_1_isBranch <= memWire_isBranch;
				memStage_1_isJAL <= memWire_isJAL;
				memStage_1_isJALR <= memWire_isJALR;
				memStage_1_isLUI <= memWire_isLUI;
				memStage_1_isAUIPC <= memWire_isAUIPC;
				memStage_1_isFence <= memWire_isFence;
				memStage_1_isSystem <= memWire_isSystem;
				memStage_1_aluOp <= memWire_aluOp;
				memStage_1_imm <= memWire_imm;
				memStage_1_rs1 <= memWire_rs1;
				memStage_1_rs2 <= memWire_rs2;
				memStage_1_rd <= memWire_rd;
				memStage_1_rs1Data <= memWire_rs1Data;
				memStage_1_rs2Data <= memWire_rs2Data;
				memStage_1_memAddr <= memWire_memAddr;
				memStage_1_memWdata <= memWire_memWdata;
				memStage_1_memRdata <= memWire_memRdata;
				memStage_1_aluResult <= memWire_aluResult;
			end
			if (_GEN_70) begin
				pcRegs_2 <= _pcRegs_T_1;
				ifStage_2_threadId <= ifWire_threadId;
				ifStage_2_pc <= ifWire_pc;
				ifStage_2_instr <= ifWire_instr;
				decStage_2_threadId <= decWire_threadId;
				decStage_2_valid <= decWire_valid;
				decStage_2_pc <= decWire_pc;
				decStage_2_instr <= decWire_instr;
				decStage_2_aluOp <= decWire_aluOp;
				decStage_2_imm <= decWire_imm;
				decStage_2_rs1 <= decWire_rs1;
				decStage_2_rs2 <= decWire_rs2;
				decStage_2_rd <= decWire_rd;
				decStage_2_rs1Data <= decWire_rs1Data;
				decStage_2_rs2Data <= decWire_rs2Data;
				decStage_2_memAddr <= decWire_memAddr;
				decStage_2_memWdata <= decWire_memWdata;
				decStage_2_memRdata <= decWire_memRdata;
				decStage_2_aluResult <= decWire_aluResult;
				exStage_2_threadId <= exWire_threadId;
				exStage_2_valid <= exWire_valid;
				exStage_2_pc <= exWire_pc;
				exStage_2_instr <= exWire_instr;
				exStage_2_isALU <= exWire_isALU;
				exStage_2_isLoad <= exWire_isLoad;
				exStage_2_isStore <= exWire_isStore;
				exStage_2_isBranch <= exWire_isBranch;
				exStage_2_isJAL <= exWire_isJAL;
				exStage_2_isJALR <= exWire_isJALR;
				exStage_2_isLUI <= exWire_isLUI;
				exStage_2_isAUIPC <= exWire_isAUIPC;
				exStage_2_isFence <= exWire_isFence;
				exStage_2_isSystem <= exWire_isSystem;
				exStage_2_aluOp <= exWire_aluOp;
				exStage_2_imm <= exWire_imm;
				exStage_2_rs1 <= exWire_rs1;
				exStage_2_rs2 <= exWire_rs2;
				exStage_2_rd <= exWire_rd;
				exStage_2_rs1Data <= exWire_rs1Data;
				exStage_2_rs2Data <= exWire_rs2Data;
				exStage_2_memAddr <= exWire_memAddr;
				exStage_2_memWdata <= exWire_memWdata;
				exStage_2_memRdata <= exWire_memRdata;
				exStage_2_aluResult <= exWire_aluResult;
				memStage_2_threadId <= memWire_threadId;
				memStage_2_valid <= memWire_valid;
				memStage_2_pc <= memWire_pc;
				memStage_2_instr <= memWire_instr;
				memStage_2_isALU <= memWire_isALU;
				memStage_2_isLoad <= memWire_isLoad;
				memStage_2_isStore <= memWire_isStore;
				memStage_2_isBranch <= memWire_isBranch;
				memStage_2_isJAL <= memWire_isJAL;
				memStage_2_isJALR <= memWire_isJALR;
				memStage_2_isLUI <= memWire_isLUI;
				memStage_2_isAUIPC <= memWire_isAUIPC;
				memStage_2_isFence <= memWire_isFence;
				memStage_2_isSystem <= memWire_isSystem;
				memStage_2_aluOp <= memWire_aluOp;
				memStage_2_imm <= memWire_imm;
				memStage_2_rs1 <= memWire_rs1;
				memStage_2_rs2 <= memWire_rs2;
				memStage_2_rd <= memWire_rd;
				memStage_2_rs1Data <= memWire_rs1Data;
				memStage_2_rs2Data <= memWire_rs2Data;
				memStage_2_memAddr <= memWire_memAddr;
				memStage_2_memWdata <= memWire_memWdata;
				memStage_2_memRdata <= memWire_memRdata;
				memStage_2_aluResult <= memWire_aluResult;
			end
			if (&currentThread) begin
				pcRegs_3 <= _pcRegs_T_1;
				ifStage_3_threadId <= ifWire_threadId;
				ifStage_3_pc <= ifWire_pc;
				ifStage_3_instr <= ifWire_instr;
				decStage_3_threadId <= decWire_threadId;
				decStage_3_valid <= decWire_valid;
				decStage_3_pc <= decWire_pc;
				decStage_3_instr <= decWire_instr;
				decStage_3_aluOp <= decWire_aluOp;
				decStage_3_imm <= decWire_imm;
				decStage_3_rs1 <= decWire_rs1;
				decStage_3_rs2 <= decWire_rs2;
				decStage_3_rd <= decWire_rd;
				decStage_3_rs1Data <= decWire_rs1Data;
				decStage_3_rs2Data <= decWire_rs2Data;
				decStage_3_memAddr <= decWire_memAddr;
				decStage_3_memWdata <= decWire_memWdata;
				decStage_3_memRdata <= decWire_memRdata;
				decStage_3_aluResult <= decWire_aluResult;
				exStage_3_threadId <= exWire_threadId;
				exStage_3_valid <= exWire_valid;
				exStage_3_pc <= exWire_pc;
				exStage_3_instr <= exWire_instr;
				exStage_3_isALU <= exWire_isALU;
				exStage_3_isLoad <= exWire_isLoad;
				exStage_3_isStore <= exWire_isStore;
				exStage_3_isBranch <= exWire_isBranch;
				exStage_3_isJAL <= exWire_isJAL;
				exStage_3_isJALR <= exWire_isJALR;
				exStage_3_isLUI <= exWire_isLUI;
				exStage_3_isAUIPC <= exWire_isAUIPC;
				exStage_3_isFence <= exWire_isFence;
				exStage_3_isSystem <= exWire_isSystem;
				exStage_3_aluOp <= exWire_aluOp;
				exStage_3_imm <= exWire_imm;
				exStage_3_rs1 <= exWire_rs1;
				exStage_3_rs2 <= exWire_rs2;
				exStage_3_rd <= exWire_rd;
				exStage_3_rs1Data <= exWire_rs1Data;
				exStage_3_rs2Data <= exWire_rs2Data;
				exStage_3_memAddr <= exWire_memAddr;
				exStage_3_memWdata <= exWire_memWdata;
				exStage_3_memRdata <= exWire_memRdata;
				exStage_3_aluResult <= exWire_aluResult;
				memStage_3_threadId <= memWire_threadId;
				memStage_3_valid <= memWire_valid;
				memStage_3_pc <= memWire_pc;
				memStage_3_instr <= memWire_instr;
				memStage_3_isALU <= memWire_isALU;
				memStage_3_isLoad <= memWire_isLoad;
				memStage_3_isStore <= memWire_isStore;
				memStage_3_isBranch <= memWire_isBranch;
				memStage_3_isJAL <= memWire_isJAL;
				memStage_3_isJALR <= memWire_isJALR;
				memStage_3_isLUI <= memWire_isLUI;
				memStage_3_isAUIPC <= memWire_isAUIPC;
				memStage_3_isFence <= memWire_isFence;
				memStage_3_isSystem <= memWire_isSystem;
				memStage_3_aluOp <= memWire_aluOp;
				memStage_3_imm <= memWire_imm;
				memStage_3_rs1 <= memWire_rs1;
				memStage_3_rs2 <= memWire_rs2;
				memStage_3_rd <= memWire_rd;
				memStage_3_rs1Data <= memWire_rs1Data;
				memStage_3_rs2Data <= memWire_rs2Data;
				memStage_3_memAddr <= memWire_memAddr;
				memStage_3_memWdata <= memWire_memWdata;
				memStage_3_memRdata <= memWire_memRdata;
				memStage_3_aluResult <= memWire_aluResult;
			end
			ifStage_0_valid <= _GEN_68 | ifStage_0_valid;
			ifStage_1_valid <= _GEN_69 | ifStage_1_valid;
			ifStage_2_valid <= _GEN_70 | ifStage_2_valid;
			ifStage_3_valid <= &currentThread | ifStage_3_valid;
			decStage_0_isALU <= (_GEN_68 ? decWire_isALU : ~_GEN_68 & decStage_0_isALU);
			decStage_0_isLoad <= (_GEN_68 ? decWire_isLoad : ~_GEN_68 & decStage_0_isLoad);
			decStage_0_isStore <= (_GEN_68 ? decWire_isStore : ~_GEN_68 & decStage_0_isStore);
			decStage_0_isBranch <= (_GEN_68 ? decWire_isBranch : ~_GEN_68 & decStage_0_isBranch);
			decStage_0_isJAL <= (_GEN_68 ? decWire_isJAL : ~_GEN_68 & decStage_0_isJAL);
			decStage_0_isJALR <= (_GEN_68 ? decWire_isJALR : ~_GEN_68 & decStage_0_isJALR);
			decStage_0_isLUI <= (_GEN_68 ? decWire_isLUI : ~_GEN_68 & decStage_0_isLUI);
			decStage_0_isAUIPC <= (_GEN_68 ? decWire_isAUIPC : ~_GEN_68 & decStage_0_isAUIPC);
			decStage_0_isFence <= (_GEN_68 ? decWire_isFence : ~_GEN_68 & decStage_0_isFence);
			decStage_0_isSystem <= (_GEN_68 ? decWire_isSystem : ~_GEN_68 & decStage_0_isSystem);
			decStage_1_isALU <= (_GEN_69 ? decWire_isALU : ~_GEN_69 & decStage_1_isALU);
			decStage_1_isLoad <= (_GEN_69 ? decWire_isLoad : ~_GEN_69 & decStage_1_isLoad);
			decStage_1_isStore <= (_GEN_69 ? decWire_isStore : ~_GEN_69 & decStage_1_isStore);
			decStage_1_isBranch <= (_GEN_69 ? decWire_isBranch : ~_GEN_69 & decStage_1_isBranch);
			decStage_1_isJAL <= (_GEN_69 ? decWire_isJAL : ~_GEN_69 & decStage_1_isJAL);
			decStage_1_isJALR <= (_GEN_69 ? decWire_isJALR : ~_GEN_69 & decStage_1_isJALR);
			decStage_1_isLUI <= (_GEN_69 ? decWire_isLUI : ~_GEN_69 & decStage_1_isLUI);
			decStage_1_isAUIPC <= (_GEN_69 ? decWire_isAUIPC : ~_GEN_69 & decStage_1_isAUIPC);
			decStage_1_isFence <= (_GEN_69 ? decWire_isFence : ~_GEN_69 & decStage_1_isFence);
			decStage_1_isSystem <= (_GEN_69 ? decWire_isSystem : ~_GEN_69 & decStage_1_isSystem);
			decStage_2_isALU <= (_GEN_70 ? decWire_isALU : ~_GEN_70 & decStage_2_isALU);
			decStage_2_isLoad <= (_GEN_70 ? decWire_isLoad : ~_GEN_70 & decStage_2_isLoad);
			decStage_2_isStore <= (_GEN_70 ? decWire_isStore : ~_GEN_70 & decStage_2_isStore);
			decStage_2_isBranch <= (_GEN_70 ? decWire_isBranch : ~_GEN_70 & decStage_2_isBranch);
			decStage_2_isJAL <= (_GEN_70 ? decWire_isJAL : ~_GEN_70 & decStage_2_isJAL);
			decStage_2_isJALR <= (_GEN_70 ? decWire_isJALR : ~_GEN_70 & decStage_2_isJALR);
			decStage_2_isLUI <= (_GEN_70 ? decWire_isLUI : ~_GEN_70 & decStage_2_isLUI);
			decStage_2_isAUIPC <= (_GEN_70 ? decWire_isAUIPC : ~_GEN_70 & decStage_2_isAUIPC);
			decStage_2_isFence <= (_GEN_70 ? decWire_isFence : ~_GEN_70 & decStage_2_isFence);
			decStage_2_isSystem <= (_GEN_70 ? decWire_isSystem : ~_GEN_70 & decStage_2_isSystem);
			decStage_3_isALU <= (&currentThread ? decWire_isALU : ~(&currentThread) & decStage_3_isALU);
			decStage_3_isLoad <= (&currentThread ? decWire_isLoad : ~(&currentThread) & decStage_3_isLoad);
			decStage_3_isStore <= (&currentThread ? decWire_isStore : ~(&currentThread) & decStage_3_isStore);
			decStage_3_isBranch <= (&currentThread ? decWire_isBranch : ~(&currentThread) & decStage_3_isBranch);
			decStage_3_isJAL <= (&currentThread ? decWire_isJAL : ~(&currentThread) & decStage_3_isJAL);
			decStage_3_isJALR <= (&currentThread ? decWire_isJALR : ~(&currentThread) & decStage_3_isJALR);
			decStage_3_isLUI <= (&currentThread ? decWire_isLUI : ~(&currentThread) & decStage_3_isLUI);
			decStage_3_isAUIPC <= (&currentThread ? decWire_isAUIPC : ~(&currentThread) & decStage_3_isAUIPC);
			decStage_3_isFence <= (&currentThread ? decWire_isFence : ~(&currentThread) & decStage_3_isFence);
			decStage_3_isSystem <= (&currentThread ? decWire_isSystem : ~(&currentThread) & decStage_3_isSystem);
		end
	initial begin : sv2v_autoblock_2
		reg [31:0] _RANDOM [0:164];
	end
	instrMem_1024x32 instrMem_ext(
		.R0_addr(_ifWire_instr_T_1),
		.R0_en(1'h1),
		.R0_clk(clock),
		.R0_data(ifWire_instr),
		.W0_addr(io_instrWriteAddr_0),
		.W0_en(io_instrWriteEnable_0),
		.W0_clk(clock),
		.W0_data(io_instrWriteData_0)
	);
	RegFileMT2R1WVec regFile(
		.clock(clock),
		.reset(reset),
		.io_threadID(currentThread),
		.io_src1(decWire_rs1),
		.io_src2(decWire_rs2),
		.io_dst1(memWire_rd),
		.io_wen(_regFile_io_wen_T_3),
		.io_dst1data(wbData),
		.io_src1data(decWire_rs1Data),
		.io_src2data(decWire_rs2Data)
	);
	TetraNyteCore_Anon alu(
		.io_a(exWire_rs1Data),
		.io_b(exWire_rs2Data),
		.io_fn(exWire_aluOp),
		.io_out(exWire_aluResult)
	);
	assign io_memAddr = io_memAddr_0;
	assign io_memWdata = io_memWdata_0;
	assign io_memWe = io_memWe_0;
endmodule
